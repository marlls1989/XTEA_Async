module xtea(in_enc_t, in_enc_f, in_enc_ack, out_enc_t, out_enc_f, out_enc_ack, key_t, key_f, key_ack, clk, reset);
input  clk, reset;
drwire add_76_21_n_1002 ();
drwire add_76_21_n_1003 ();
drwire add_76_21_n_1004 ();
drwire add_76_21_n_1005 ();
drwire add_76_21_n_1006 ();
drwire add_76_21_n_1009 ();
drwire add_76_21_n_1010 ();
drwire add_76_21_n_1011 ();
drwire add_76_21_n_1012 ();
drwire add_76_21_n_1014 ();
drwire add_76_21_n_1015 ();
drwire add_76_21_n_1016 ();
drwire add_76_21_n_1017 ();
drwire add_76_21_n_1018 ();
drwire add_76_21_n_1019 ();
drwire add_76_21_n_1020 ();
drwire add_76_21_n_1031 ();
drwire add_76_21_n_1032 ();
drwire add_76_21_n_1033 ();
drwire add_76_21_n_1034 ();
drwire add_76_21_n_1035 ();
drwire add_76_21_n_1038 ();
drwire add_76_21_n_1039 ();
drwire add_76_21_n_1040 ();
drwire add_76_21_n_1041 ();
drwire add_76_21_n_1042 ();
drwire add_76_21_n_1043 ();
drwire add_76_21_n_1044 ();
drwire add_76_21_n_1045 ();
drwire add_76_21_n_1047 ();
drwire add_76_21_n_1052 ();
drwire add_76_21_n_1055 ();
drwire add_76_21_n_1056 ();
drwire add_76_21_n_1057 ();
drwire add_76_21_n_1058 ();
drwire add_76_21_n_1059 ();
drwire add_76_21_n_1060 ();
drwire add_76_21_n_1062 ();
drwire add_76_21_n_1063 ();
drwire add_76_21_n_1064 ();
drwire add_76_21_n_1065 ();
drwire add_76_21_n_1067 ();
drwire add_76_21_n_1068 ();
drwire add_76_21_n_1069 ();
drwire add_76_21_n_1070 ();
drwire add_76_21_n_1071 ();
drwire add_76_21_n_1072 ();
drwire add_76_21_n_1073 ();
drwire add_76_21_n_1074 ();
drwire add_76_21_n_1075 ();
drwire add_76_21_n_1078 ();
drwire add_76_21_n_1080 ();
drwire add_76_21_n_1082 ();
drwire add_76_21_n_1083 ();
drwire add_76_21_n_1085 ();
drwire add_76_21_n_1086 ();
drwire add_76_21_n_1088 ();
drwire add_76_21_n_1093 ();
drwire add_76_21_n_1117 ();
drwire add_76_21_n_1119 ();
drwire add_76_21_n_1121 ();
drwire add_76_21_n_1122 ();
drwire add_76_21_n_1124 ();
drwire add_76_21_n_1127 ();
drwire add_76_21_n_1130 ();
drwire add_76_21_n_1134 ();
drwire add_76_21_n_1135 ();
drwire add_76_21_n_1137 ();
drwire add_76_21_n_1141 ();
drwire add_76_21_n_1144 ();
drwire add_76_21_n_1148 ();
drwire add_76_21_n_1150 ();
drwire add_76_21_n_1155 ();
drwire add_76_21_n_1156 ();
drwire add_76_21_n_1158 ();
drwire add_76_21_n_1160 ();
drwire add_76_21_n_1161 ();
drwire add_76_21_n_1163 ();
drwire add_76_21_n_1165 ();
drwire add_76_21_n_1167 ();
drwire add_76_21_n_1170 ();
drwire add_76_21_n_1172 ();
drwire add_76_21_n_1173 ();
drwire add_76_21_n_1174 ();
drwire add_76_21_n_1176 ();
drwire add_76_21_n_1178 ();
drwire add_76_21_n_1181 ();
drwire add_76_21_n_1183 ();
drwire add_76_21_n_1185 ();
drwire add_76_21_n_1192 ();
drwire add_76_21_n_1194 ();
drwire add_76_21_n_1195 ();
drwire add_76_21_n_1200 ();
drwire add_76_21_n_1203 ();
drwire add_76_21_n_1207 ();
drwire add_76_21_n_1209 ();
drwire add_76_21_n_1216 ();
drwire add_76_21_n_1230 ();
drwire add_76_21_n_1231 ();
drwire add_76_21_n_1233 ();
drwire add_76_21_n_1235 ();
drwire add_76_21_n_1237 ();
drwire add_76_21_n_1238 ();
drwire add_76_21_n_1240 ();
drwire add_76_21_n_1242 ();
drwire add_76_21_n_1244 ();
drwire add_76_21_n_1249 ();
drwire add_76_21_n_1251 ();
drwire add_76_21_n_1254 ();
drwire add_76_21_n_1256 ();
drwire add_76_21_n_1261 ();
drwire add_76_21_n_1263 ();
drwire add_76_21_n_1267 ();
drwire add_76_21_n_1272 ();
drwire add_76_21_n_1274 ();
drwire add_76_21_n_1277 ();
drwire add_76_21_n_1394 ();
drwire add_76_21_n_1395 ();
drwire add_76_21_n_799 ();
drwire add_76_21_n_800 ();
drwire add_76_21_n_804 ();
drwire add_76_21_n_805 ();
drwire add_76_21_n_811 ();
drwire add_76_21_n_815 ();
drwire add_76_21_n_817 ();
drwire add_76_21_n_818 ();
drwire add_76_21_n_819 ();
drwire add_76_21_n_820 ();
drwire add_76_21_n_824 ();
drwire add_76_21_n_835 ();
drwire add_76_21_n_837 ();
drwire add_76_21_n_846 ();
drwire add_76_21_n_851 ();
drwire add_76_21_n_854 ();
drwire add_76_21_n_858 ();
drwire add_76_21_n_859 ();
drwire add_76_21_n_861 ();
drwire add_76_21_n_863 ();
drwire add_76_21_n_872 ();
drwire add_76_21_n_875 ();
drwire add_76_21_n_878 ();
drwire add_76_21_n_881 ();
drwire add_76_21_n_882 ();
drwire add_76_21_n_884 ();
drwire add_76_21_n_886 ();
drwire add_76_21_n_888 ();
drwire add_76_21_n_889 ();
drwire add_76_21_n_890 ();
drwire add_76_21_n_891 ();
drwire add_76_21_n_893 ();
drwire add_76_21_n_894 ();
drwire add_76_21_n_896 ();
drwire add_76_21_n_900 ();
drwire add_76_21_n_902 ();
drwire add_76_21_n_905 ();
drwire add_76_21_n_906 ();
drwire add_76_21_n_907 ();
drwire add_76_21_n_908 ();
drwire add_76_21_n_911 ();
drwire add_76_21_n_912 ();
drwire add_76_21_n_913 ();
drwire add_76_21_n_914 ();
drwire add_76_21_n_915 ();
drwire add_76_21_n_918 ();
drwire add_76_21_n_919 ();
drwire add_76_21_n_922 ();
drwire add_76_21_n_925 ();
drwire add_76_21_n_926 ();
drwire add_76_21_n_928 ();
drwire add_76_21_n_929 ();
drwire add_76_21_n_930 ();
drwire add_76_21_n_932 ();
drwire add_76_21_n_935 ();
drwire add_76_21_n_936 ();
drwire add_76_21_n_938 ();
drwire add_76_21_n_940 ();
drwire add_76_21_n_942 ();
drwire add_76_21_n_947 ();
drwire add_76_21_n_948 ();
drwire add_76_21_n_949 ();
drwire add_76_21_n_950 ();
drwire add_76_21_n_951 ();
drwire add_76_21_n_957 ();
drwire add_76_21_n_959 ();
drwire add_76_21_n_961 ();
drwire add_76_21_n_963 ();
drwire add_76_21_n_964 ();
drwire add_76_21_n_966 ();
drwire add_76_21_n_968 ();
drwire add_76_21_n_971 ();
drwire add_76_21_n_975 ();
drwire add_76_21_n_977 ();
drwire add_76_21_n_978 ();
drwire add_76_21_n_980 ();
drwire add_76_21_n_981 ();
drwire add_76_21_n_982 ();
drwire add_76_21_n_984 ();
drwire add_76_21_n_985 ();
drwire add_76_21_n_988 ();
drwire add_76_21_n_990 ();
drwire add_76_21_n_992 ();
drwire add_76_21_n_995 ();
drwire add_76_69_n_1000 ();
drwire add_76_69_n_1001 ();
drwire add_76_69_n_1002 ();
drwire add_76_69_n_1003 ();
drwire add_76_69_n_1004 ();
drwire add_76_69_n_1005 ();
drwire add_76_69_n_1006 ();
drwire add_76_69_n_1007 ();
drwire add_76_69_n_1008 ();
drwire add_76_69_n_1009 ();
drwire add_76_69_n_1010 ();
drwire add_76_69_n_1011 ();
drwire add_76_69_n_1012 ();
drwire add_76_69_n_1013 ();
drwire add_76_69_n_1014 ();
drwire add_76_69_n_1015 ();
drwire add_76_69_n_1016 ();
drwire add_76_69_n_1017 ();
drwire add_76_69_n_1018 ();
drwire add_76_69_n_1019 ();
drwire add_76_69_n_1020 ();
drwire add_76_69_n_1021 ();
drwire add_76_69_n_1022 ();
drwire add_76_69_n_1023 ();
drwire add_76_69_n_1024 ();
drwire add_76_69_n_1025 ();
drwire add_76_69_n_1026 ();
drwire add_76_69_n_1027 ();
drwire add_76_69_n_1028 ();
drwire add_76_69_n_1029 ();
drwire add_76_69_n_1030 ();
drwire add_76_69_n_1031 ();
drwire add_76_69_n_1032 ();
drwire add_76_69_n_1033 ();
drwire add_76_69_n_1034 ();
drwire add_76_69_n_1035 ();
drwire add_76_69_n_1036 ();
drwire add_76_69_n_1037 ();
drwire add_76_69_n_1038 ();
drwire add_76_69_n_1039 ();
drwire add_76_69_n_1040 ();
drwire add_76_69_n_1041 ();
drwire add_76_69_n_1042 ();
drwire add_76_69_n_1043 ();
drwire add_76_69_n_1044 ();
drwire add_76_69_n_1046 ();
drwire add_76_69_n_1047 ();
drwire add_76_69_n_1048 ();
drwire add_76_69_n_1051 ();
drwire add_76_69_n_1060 ();
drwire add_76_69_n_1066 ();
drwire add_76_69_n_1067 ();
drwire add_76_69_n_1068 ();
drwire add_76_69_n_1069 ();
drwire add_76_69_n_1070 ();
drwire add_76_69_n_1071 ();
drwire add_76_69_n_1072 ();
drwire add_76_69_n_1073 ();
drwire add_76_69_n_1074 ();
drwire add_76_69_n_1075 ();
drwire add_76_69_n_1076 ();
drwire add_76_69_n_1077 ();
drwire add_76_69_n_1078 ();
drwire add_76_69_n_1079 ();
drwire add_76_69_n_1080 ();
drwire add_76_69_n_1081 ();
drwire add_76_69_n_1082 ();
drwire add_76_69_n_1083 ();
drwire add_76_69_n_1084 ();
drwire add_76_69_n_1085 ();
drwire add_76_69_n_1086 ();
drwire add_76_69_n_1087 ();
drwire add_76_69_n_1088 ();
drwire add_76_69_n_1090 ();
drwire add_76_69_n_1091 ();
drwire add_76_69_n_1092 ();
drwire add_76_69_n_1093 ();
drwire add_76_69_n_1094 ();
drwire add_76_69_n_1095 ();
drwire add_76_69_n_1096 ();
drwire add_76_69_n_1097 ();
drwire add_76_69_n_1098 ();
drwire add_76_69_n_1099 ();
drwire add_76_69_n_1100 ();
drwire add_76_69_n_1101 ();
drwire add_76_69_n_1102 ();
drwire add_76_69_n_1103 ();
drwire add_76_69_n_1104 ();
drwire add_76_69_n_1105 ();
drwire add_76_69_n_1106 ();
drwire add_76_69_n_1107 ();
drwire add_76_69_n_1108 ();
drwire add_76_69_n_1109 ();
drwire add_76_69_n_1110 ();
drwire add_76_69_n_1111 ();
drwire add_76_69_n_1114 ();
drwire add_76_69_n_1117 ();
drwire add_76_69_n_1119 ();
drwire add_76_69_n_625 ();
drwire add_76_69_n_631 ();
drwire add_76_69_n_651 ();
drwire add_76_69_n_653 ();
drwire add_76_69_n_654 ();
drwire add_76_69_n_655 ();
drwire add_76_69_n_656 ();
drwire add_76_69_n_658 ();
drwire add_76_69_n_659 ();
drwire add_76_69_n_660 ();
drwire add_76_69_n_661 ();
drwire add_76_69_n_664 ();
drwire add_76_69_n_665 ();
drwire add_76_69_n_666 ();
drwire add_76_69_n_668 ();
drwire add_76_69_n_669 ();
drwire add_76_69_n_674 ();
drwire add_76_69_n_683 ();
drwire add_76_69_n_684 ();
drwire add_76_69_n_685 ();
drwire add_76_69_n_690 ();
drwire add_76_69_n_692 ();
drwire add_76_69_n_696 ();
drwire add_76_69_n_697 ();
drwire add_76_69_n_698 ();
drwire add_76_69_n_699 ();
drwire add_76_69_n_700 ();
drwire add_76_69_n_701 ();
drwire add_76_69_n_705 ();
drwire add_76_69_n_706 ();
drwire add_76_69_n_707 ();
drwire add_76_69_n_709 ();
drwire add_76_69_n_710 ();
drwire add_76_69_n_711 ();
drwire add_76_69_n_714 ();
drwire add_76_69_n_715 ();
drwire add_76_69_n_716 ();
drwire add_76_69_n_717 ();
drwire add_76_69_n_722 ();
drwire add_76_69_n_723 ();
drwire add_76_69_n_727 ();
drwire add_76_69_n_729 ();
drwire add_76_69_n_732 ();
drwire add_76_69_n_734 ();
drwire add_76_69_n_735 ();
drwire add_76_69_n_736 ();
drwire add_76_69_n_737 ();
drwire add_76_69_n_738 ();
drwire add_76_69_n_740 ();
drwire add_76_69_n_741 ();
drwire add_76_69_n_742 ();
drwire add_76_69_n_743 ();
drwire add_76_69_n_744 ();
drwire add_76_69_n_745 ();
drwire add_76_69_n_746 ();
drwire add_76_69_n_748 ();
drwire add_76_69_n_749 ();
drwire add_76_69_n_750 ();
drwire add_76_69_n_753 ();
drwire add_76_69_n_755 ();
drwire add_76_69_n_756 ();
drwire add_76_69_n_757 ();
drwire add_76_69_n_759 ();
drwire add_76_69_n_760 ();
drwire add_76_69_n_761 ();
drwire add_76_69_n_762 ();
drwire add_76_69_n_763 ();
drwire add_76_69_n_765 ();
drwire add_76_69_n_766 ();
drwire add_76_69_n_767 ();
drwire add_76_69_n_768 ();
drwire add_76_69_n_771 ();
drwire add_76_69_n_772 ();
drwire add_76_69_n_774 ();
drwire add_76_69_n_776 ();
drwire add_76_69_n_778 ();
drwire add_76_69_n_779 ();
drwire add_76_69_n_780 ();
drwire add_76_69_n_781 ();
drwire add_76_69_n_782 ();
drwire add_76_69_n_783 ();
drwire add_76_69_n_786 ();
drwire add_76_69_n_788 ();
drwire add_76_69_n_791 ();
drwire add_76_69_n_793 ();
drwire add_76_69_n_794 ();
drwire add_76_69_n_795 ();
drwire add_76_69_n_797 ();
drwire add_76_69_n_799 ();
drwire add_76_69_n_800 ();
drwire add_76_69_n_802 ();
drwire add_76_69_n_806 ();
drwire add_76_69_n_807 ();
drwire add_76_69_n_809 ();
drwire add_76_69_n_810 ();
drwire add_76_69_n_812 ();
drwire add_76_69_n_813 ();
drwire add_76_69_n_815 ();
drwire add_76_69_n_819 ();
drwire add_76_69_n_820 ();
drwire add_76_69_n_821 ();
drwire add_76_69_n_823 ();
drwire add_76_69_n_825 ();
drwire add_76_69_n_831 ();
drwire add_76_69_n_832 ();
drwire add_76_69_n_833 ();
drwire add_76_69_n_834 ();
drwire add_76_69_n_835 ();
drwire add_76_69_n_836 ();
drwire add_76_69_n_837 ();
drwire add_76_69_n_838 ();
drwire add_76_69_n_839 ();
drwire add_76_69_n_840 ();
drwire add_76_69_n_841 ();
drwire add_76_69_n_842 ();
drwire add_76_69_n_843 ();
drwire add_76_69_n_844 ();
drwire add_76_69_n_845 ();
drwire add_76_69_n_846 ();
drwire add_76_69_n_847 ();
drwire add_76_69_n_851 ();
drwire add_76_69_n_852 ();
drwire add_76_69_n_860 ();
drwire add_76_69_n_861 ();
drwire add_76_69_n_862 ();
drwire add_76_69_n_863 ();
drwire add_76_69_n_864 ();
drwire add_76_69_n_867 ();
drwire add_76_69_n_868 ();
drwire add_76_69_n_869 ();
drwire add_76_69_n_870 ();
drwire add_76_69_n_872 ();
drwire add_76_69_n_874 ();
drwire add_76_69_n_875 ();
drwire add_76_69_n_877 ();
drwire add_76_69_n_878 ();
drwire add_76_69_n_879 ();
drwire add_76_69_n_883 ();
drwire add_76_69_n_884 ();
drwire add_76_69_n_885 ();
drwire add_76_69_n_886 ();
drwire add_76_69_n_887 ();
drwire add_76_69_n_888 ();
drwire add_76_69_n_889 ();
drwire add_76_69_n_890 ();
drwire add_76_69_n_893 ();
drwire add_76_69_n_894 ();
drwire add_76_69_n_895 ();
drwire add_76_69_n_896 ();
drwire add_76_69_n_897 ();
drwire add_76_69_n_898 ();
drwire add_76_69_n_899 ();
drwire add_76_69_n_900 ();
drwire add_76_69_n_901 ();
drwire add_76_69_n_902 ();
drwire add_76_69_n_903 ();
drwire add_76_69_n_905 ();
drwire add_76_69_n_907 ();
drwire add_76_69_n_908 ();
drwire add_76_69_n_909 ();
drwire add_76_69_n_911 ();
drwire add_76_69_n_912 ();
drwire add_76_69_n_913 ();
drwire add_76_69_n_915 ();
drwire add_76_69_n_918 ();
drwire add_76_69_n_919 ();
drwire add_76_69_n_921 ();
drwire add_76_69_n_923 ();
drwire add_76_69_n_925 ();
drwire add_76_69_n_927 ();
drwire add_76_69_n_935 ();
drwire add_76_69_n_948 ();
drwire add_76_69_n_952 ();
drwire add_76_69_n_954 ();
drwire add_76_69_n_964 ();
drwire add_76_69_n_977 ();
drwire add_76_69_n_981 ();
drwire add_76_69_n_983 ();
drwire add_76_69_n_988 ();
drwire add_76_69_n_994 ();
drwire add_76_69_n_995 ();
drwire add_76_69_n_997 ();
drwire add_76_69_n_998 ();
drwire add_76_69_n_999 ();
drwire add_76_82_n_1000 ();
drwire add_76_82_n_1004 ();
drwire add_76_82_n_1005 ();
drwire add_76_82_n_1007 ();
drwire add_76_82_n_1009 ();
drwire add_76_82_n_1010 ();
drwire add_76_82_n_1012 ();
drwire add_76_82_n_1013 ();
drwire add_76_82_n_1015 ();
drwire add_76_82_n_1018 ();
drwire add_76_82_n_1019 ();
drwire add_76_82_n_1020 ();
drwire add_76_82_n_1022 ();
drwire add_76_82_n_1028 ();
drwire add_76_82_n_1030 ();
drwire add_76_82_n_1031 ();
drwire add_76_82_n_1032 ();
drwire add_76_82_n_1034 ();
drwire add_76_82_n_1035 ();
drwire add_76_82_n_1036 ();
drwire add_76_82_n_1037 ();
drwire add_76_82_n_1038 ();
drwire add_76_82_n_1039 ();
drwire add_76_82_n_1040 ();
drwire add_76_82_n_1041 ();
drwire add_76_82_n_1042 ();
drwire add_76_82_n_1044 ();
drwire add_76_82_n_1048 ();
drwire add_76_82_n_1049 ();
drwire add_76_82_n_1057 ();
drwire add_76_82_n_1058 ();
drwire add_76_82_n_1059 ();
drwire add_76_82_n_1060 ();
drwire add_76_82_n_1061 ();
drwire add_76_82_n_1062 ();
drwire add_76_82_n_1063 ();
drwire add_76_82_n_1064 ();
drwire add_76_82_n_1066 ();
drwire add_76_82_n_1068 ();
drwire add_76_82_n_1069 ();
drwire add_76_82_n_1070 ();
drwire add_76_82_n_1072 ();
drwire add_76_82_n_1073 ();
drwire add_76_82_n_1075 ();
drwire add_76_82_n_1080 ();
drwire add_76_82_n_1081 ();
drwire add_76_82_n_1082 ();
drwire add_76_82_n_1083 ();
drwire add_76_82_n_1084 ();
drwire add_76_82_n_1085 ();
drwire add_76_82_n_1086 ();
drwire add_76_82_n_1087 ();
drwire add_76_82_n_1088 ();
drwire add_76_82_n_1089 ();
drwire add_76_82_n_1090 ();
drwire add_76_82_n_1091 ();
drwire add_76_82_n_1092 ();
drwire add_76_82_n_1093 ();
drwire add_76_82_n_1094 ();
drwire add_76_82_n_1095 ();
drwire add_76_82_n_1096 ();
drwire add_76_82_n_1097 ();
drwire add_76_82_n_1098 ();
drwire add_76_82_n_1100 ();
drwire add_76_82_n_1102 ();
drwire add_76_82_n_1104 ();
drwire add_76_82_n_1106 ();
drwire add_76_82_n_1109 ();
drwire add_76_82_n_1111 ();
drwire add_76_82_n_1112 ();
drwire add_76_82_n_1113 ();
drwire add_76_82_n_1114 ();
drwire add_76_82_n_1116 ();
drwire add_76_82_n_1117 ();
drwire add_76_82_n_1122 ();
drwire add_76_82_n_1144 ();
drwire add_76_82_n_1148 ();
drwire add_76_82_n_1153 ();
drwire add_76_82_n_1168 ();
drwire add_76_82_n_1191 ();
drwire add_76_82_n_1194 ();
drwire add_76_82_n_1196 ();
drwire add_76_82_n_1198 ();
drwire add_76_82_n_1199 ();
drwire add_76_82_n_1200 ();
drwire add_76_82_n_1201 ();
drwire add_76_82_n_1203 ();
drwire add_76_82_n_1204 ();
drwire add_76_82_n_1205 ();
drwire add_76_82_n_1206 ();
drwire add_76_82_n_1207 ();
drwire add_76_82_n_1208 ();
drwire add_76_82_n_1209 ();
drwire add_76_82_n_1210 ();
drwire add_76_82_n_1211 ();
drwire add_76_82_n_1212 ();
drwire add_76_82_n_1213 ();
drwire add_76_82_n_1214 ();
drwire add_76_82_n_1215 ();
drwire add_76_82_n_1216 ();
drwire add_76_82_n_1217 ();
drwire add_76_82_n_1218 ();
drwire add_76_82_n_1219 ();
drwire add_76_82_n_1222 ();
drwire add_76_82_n_1223 ();
drwire add_76_82_n_1224 ();
drwire add_76_82_n_1225 ();
drwire add_76_82_n_1226 ();
drwire add_76_82_n_1227 ();
drwire add_76_82_n_1228 ();
drwire add_76_82_n_1229 ();
drwire add_76_82_n_1230 ();
drwire add_76_82_n_1231 ();
drwire add_76_82_n_1232 ();
drwire add_76_82_n_1233 ();
drwire add_76_82_n_1234 ();
drwire add_76_82_n_1235 ();
drwire add_76_82_n_1236 ();
drwire add_76_82_n_1237 ();
drwire add_76_82_n_1238 ();
drwire add_76_82_n_1239 ();
drwire add_76_82_n_1242 ();
drwire add_76_82_n_1243 ();
drwire add_76_82_n_1257 ();
drwire add_76_82_n_1258 ();
drwire add_76_82_n_1259 ();
drwire add_76_82_n_1260 ();
drwire add_76_82_n_1261 ();
drwire add_76_82_n_1262 ();
drwire add_76_82_n_1263 ();
drwire add_76_82_n_1264 ();
drwire add_76_82_n_1265 ();
drwire add_76_82_n_1266 ();
drwire add_76_82_n_1267 ();
drwire add_76_82_n_1268 ();
drwire add_76_82_n_1269 ();
drwire add_76_82_n_1270 ();
drwire add_76_82_n_1271 ();
drwire add_76_82_n_1272 ();
drwire add_76_82_n_1273 ();
drwire add_76_82_n_1274 ();
drwire add_76_82_n_1275 ();
drwire add_76_82_n_1276 ();
drwire add_76_82_n_1277 ();
drwire add_76_82_n_1278 ();
drwire add_76_82_n_1279 ();
drwire add_76_82_n_1284 ();
drwire add_76_82_n_1285 ();
drwire add_76_82_n_1286 ();
drwire add_76_82_n_1287 ();
drwire add_76_82_n_1289 ();
drwire add_76_82_n_1290 ();
drwire add_76_82_n_1291 ();
drwire add_76_82_n_1292 ();
drwire add_76_82_n_1293 ();
drwire add_76_82_n_1294 ();
drwire add_76_82_n_1295 ();
drwire add_76_82_n_1296 ();
drwire add_76_82_n_1297 ();
drwire add_76_82_n_1298 ();
drwire add_76_82_n_1299 ();
drwire add_76_82_n_1300 ();
drwire add_76_82_n_1301 ();
drwire add_76_82_n_1302 ();
drwire add_76_82_n_1303 ();
drwire add_76_82_n_1306 ();
drwire add_76_82_n_1307 ();
drwire add_76_82_n_1308 ();
drwire add_76_82_n_1311 ();
drwire add_76_82_n_1318 ();
drwire add_76_82_n_815 ();
drwire add_76_82_n_820 ();
drwire add_76_82_n_839 ();
drwire add_76_82_n_840 ();
drwire add_76_82_n_842 ();
drwire add_76_82_n_846 ();
drwire add_76_82_n_847 ();
drwire add_76_82_n_848 ();
drwire add_76_82_n_849 ();
drwire add_76_82_n_850 ();
drwire add_76_82_n_853 ();
drwire add_76_82_n_854 ();
drwire add_76_82_n_855 ();
drwire add_76_82_n_856 ();
drwire add_76_82_n_858 ();
drwire add_76_82_n_863 ();
drwire add_76_82_n_864 ();
drwire add_76_82_n_879 ();
drwire add_76_82_n_885 ();
drwire add_76_82_n_888 ();
drwire add_76_82_n_892 ();
drwire add_76_82_n_893 ();
drwire add_76_82_n_895 ();
drwire add_76_82_n_896 ();
drwire add_76_82_n_898 ();
drwire add_76_82_n_901 ();
drwire add_76_82_n_902 ();
drwire add_76_82_n_903 ();
drwire add_76_82_n_904 ();
drwire add_76_82_n_905 ();
drwire add_76_82_n_908 ();
drwire add_76_82_n_909 ();
drwire add_76_82_n_910 ();
drwire add_76_82_n_911 ();
drwire add_76_82_n_915 ();
drwire add_76_82_n_916 ();
drwire add_76_82_n_918 ();
drwire add_76_82_n_920 ();
drwire add_76_82_n_922 ();
drwire add_76_82_n_923 ();
drwire add_76_82_n_928 ();
drwire add_76_82_n_930 ();
drwire add_76_82_n_931 ();
drwire add_76_82_n_933 ();
drwire add_76_82_n_934 ();
drwire add_76_82_n_936 ();
drwire add_76_82_n_937 ();
drwire add_76_82_n_938 ();
drwire add_76_82_n_939 ();
drwire add_76_82_n_940 ();
drwire add_76_82_n_941 ();
drwire add_76_82_n_944 ();
drwire add_76_82_n_945 ();
drwire add_76_82_n_946 ();
drwire add_76_82_n_948 ();
drwire add_76_82_n_949 ();
drwire add_76_82_n_951 ();
drwire add_76_82_n_954 ();
drwire add_76_82_n_955 ();
drwire add_76_82_n_956 ();
drwire add_76_82_n_959 ();
drwire add_76_82_n_960 ();
drwire add_76_82_n_961 ();
drwire add_76_82_n_963 ();
drwire add_76_82_n_966 ();
drwire add_76_82_n_967 ();
drwire add_76_82_n_969 ();
drwire add_76_82_n_971 ();
drwire add_76_82_n_974 ();
drwire add_76_82_n_975 ();
drwire add_76_82_n_976 ();
drwire add_76_82_n_979 ();
drwire add_76_82_n_980 ();
drwire add_76_82_n_981 ();
drwire add_76_82_n_984 ();
drwire add_76_82_n_986 ();
drwire add_76_82_n_989 ();
drwire add_76_82_n_991 ();
drwire add_76_82_n_992 ();
drwire add_76_82_n_996 ();
drwire add_76_82_n_998 ();
drwire add_88_21_n_1000 ();
drwire add_88_21_n_1002 ();
drwire add_88_21_n_1003 ();
drwire add_88_21_n_1005 ();
drwire add_88_21_n_1006 ();
drwire add_88_21_n_1008 ();
drwire add_88_21_n_1010 ();
drwire add_88_21_n_1012 ();
drwire add_88_21_n_1013 ();
drwire add_88_21_n_1014 ();
drwire add_88_21_n_1015 ();
drwire add_88_21_n_1020 ();
drwire add_88_21_n_1022 ();
drwire add_88_21_n_1023 ();
drwire add_88_21_n_1024 ();
drwire add_88_21_n_1026 ();
drwire add_88_21_n_1028 ();
drwire add_88_21_n_1030 ();
drwire add_88_21_n_1032 ();
drwire add_88_21_n_1033 ();
drwire add_88_21_n_1035 ();
drwire add_88_21_n_1037 ();
drwire add_88_21_n_1039 ();
drwire add_88_21_n_1042 ();
drwire add_88_21_n_1043 ();
drwire add_88_21_n_1049 ();
drwire add_88_21_n_1050 ();
drwire add_88_21_n_1053 ();
drwire add_88_21_n_1055 ();
drwire add_88_21_n_1060 ();
drwire add_88_21_n_1062 ();
drwire add_88_21_n_1063 ();
drwire add_88_21_n_1064 ();
drwire add_88_21_n_1067 ();
drwire add_88_21_n_1072 ();
drwire add_88_21_n_1093 ();
drwire add_88_21_n_1095 ();
drwire add_88_21_n_1097 ();
drwire add_88_21_n_1098 ();
drwire add_88_21_n_1099 ();
drwire add_88_21_n_1101 ();
drwire add_88_21_n_1103 ();
drwire add_88_21_n_1105 ();
drwire add_88_21_n_1107 ();
drwire add_88_21_n_1108 ();
drwire add_88_21_n_1111 ();
drwire add_88_21_n_1112 ();
drwire add_88_21_n_1113 ();
drwire add_88_21_n_1117 ();
drwire add_88_21_n_1118 ();
drwire add_88_21_n_1119 ();
drwire add_88_21_n_1121 ();
drwire add_88_21_n_1122 ();
drwire add_88_21_n_1123 ();
drwire add_88_21_n_1126 ();
drwire add_88_21_n_1127 ();
drwire add_88_21_n_1129 ();
drwire add_88_21_n_1131 ();
drwire add_88_21_n_1132 ();
drwire add_88_21_n_1133 ();
drwire add_88_21_n_1134 ();
drwire add_88_21_n_1138 ();
drwire add_88_21_n_1139 ();
drwire add_88_21_n_1140 ();
drwire add_88_21_n_1142 ();
drwire add_88_21_n_1255 ();
drwire add_88_21_n_1256 ();
drwire add_88_21_n_673 ();
drwire add_88_21_n_681 ();
drwire add_88_21_n_688 ();
drwire add_88_21_n_693 ();
drwire add_88_21_n_713 ();
drwire add_88_21_n_715 ();
drwire add_88_21_n_716 ();
drwire add_88_21_n_718 ();
drwire add_88_21_n_720 ();
drwire add_88_21_n_721 ();
drwire add_88_21_n_726 ();
drwire add_88_21_n_727 ();
drwire add_88_21_n_731 ();
drwire add_88_21_n_733 ();
drwire add_88_21_n_734 ();
drwire add_88_21_n_735 ();
drwire add_88_21_n_741 ();
drwire add_88_21_n_742 ();
drwire add_88_21_n_743 ();
drwire add_88_21_n_744 ();
drwire add_88_21_n_746 ();
drwire add_88_21_n_747 ();
drwire add_88_21_n_749 ();
drwire add_88_21_n_750 ();
drwire add_88_21_n_751 ();
drwire add_88_21_n_753 ();
drwire add_88_21_n_756 ();
drwire add_88_21_n_758 ();
drwire add_88_21_n_760 ();
drwire add_88_21_n_762 ();
drwire add_88_21_n_764 ();
drwire add_88_21_n_768 ();
drwire add_88_21_n_769 ();
drwire add_88_21_n_771 ();
drwire add_88_21_n_772 ();
drwire add_88_21_n_773 ();
drwire add_88_21_n_774 ();
drwire add_88_21_n_775 ();
drwire add_88_21_n_778 ();
drwire add_88_21_n_779 ();
drwire add_88_21_n_780 ();
drwire add_88_21_n_781 ();
drwire add_88_21_n_783 ();
drwire add_88_21_n_787 ();
drwire add_88_21_n_788 ();
drwire add_88_21_n_789 ();
drwire add_88_21_n_791 ();
drwire add_88_21_n_793 ();
drwire add_88_21_n_795 ();
drwire add_88_21_n_796 ();
drwire add_88_21_n_797 ();
drwire add_88_21_n_799 ();
drwire add_88_21_n_800 ();
drwire add_88_21_n_801 ();
drwire add_88_21_n_803 ();
drwire add_88_21_n_805 ();
drwire add_88_21_n_806 ();
drwire add_88_21_n_810 ();
drwire add_88_21_n_812 ();
drwire add_88_21_n_813 ();
drwire add_88_21_n_815 ();
drwire add_88_21_n_819 ();
drwire add_88_21_n_820 ();
drwire add_88_21_n_823 ();
drwire add_88_21_n_825 ();
drwire add_88_21_n_826 ();
drwire add_88_21_n_828 ();
drwire add_88_21_n_830 ();
drwire add_88_21_n_833 ();
drwire add_88_21_n_834 ();
drwire add_88_21_n_838 ();
drwire add_88_21_n_839 ();
drwire add_88_21_n_840 ();
drwire add_88_21_n_841 ();
drwire add_88_21_n_843 ();
drwire add_88_21_n_845 ();
drwire add_88_21_n_847 ();
drwire add_88_21_n_848 ();
drwire add_88_21_n_850 ();
drwire add_88_21_n_852 ();
drwire add_88_21_n_856 ();
drwire add_88_21_n_857 ();
drwire add_88_21_n_859 ();
drwire add_88_21_n_860 ();
drwire add_88_21_n_865 ();
drwire add_88_21_n_866 ();
drwire add_88_21_n_868 ();
drwire add_88_21_n_869 ();
drwire add_88_21_n_870 ();
drwire add_88_21_n_871 ();
drwire add_88_21_n_872 ();
drwire add_88_21_n_873 ();
drwire add_88_21_n_874 ();
drwire add_88_21_n_875 ();
drwire add_88_21_n_876 ();
drwire add_88_21_n_877 ();
drwire add_88_21_n_878 ();
drwire add_88_21_n_882 ();
drwire add_88_21_n_883 ();
drwire add_88_21_n_884 ();
drwire add_88_21_n_887 ();
drwire add_88_21_n_895 ();
drwire add_88_21_n_896 ();
drwire add_88_21_n_897 ();
drwire add_88_21_n_898 ();
drwire add_88_21_n_899 ();
drwire add_88_21_n_900 ();
drwire add_88_21_n_901 ();
drwire add_88_21_n_902 ();
drwire add_88_21_n_903 ();
drwire add_88_21_n_904 ();
drwire add_88_21_n_905 ();
drwire add_88_21_n_906 ();
drwire add_88_21_n_907 ();
drwire add_88_21_n_909 ();
drwire add_88_21_n_910 ();
drwire add_88_21_n_911 ();
drwire add_88_21_n_913 ();
drwire add_88_21_n_914 ();
drwire add_88_21_n_915 ();
drwire add_88_21_n_916 ();
drwire add_88_21_n_917 ();
drwire add_88_21_n_918 ();
drwire add_88_21_n_919 ();
drwire add_88_21_n_920 ();
drwire add_88_21_n_921 ();
drwire add_88_21_n_923 ();
drwire add_88_21_n_924 ();
drwire add_88_21_n_925 ();
drwire add_88_21_n_926 ();
drwire add_88_21_n_927 ();
drwire add_88_21_n_928 ();
drwire add_88_21_n_929 ();
drwire add_88_21_n_930 ();
drwire add_88_21_n_931 ();
drwire add_88_21_n_933 ();
drwire add_88_21_n_934 ();
drwire add_88_21_n_935 ();
drwire add_88_21_n_937 ();
drwire add_88_21_n_939 ();
drwire add_88_21_n_941 ();
drwire add_88_21_n_942 ();
drwire add_88_21_n_944 ();
drwire add_88_21_n_946 ();
drwire add_88_21_n_947 ();
drwire add_88_21_n_949 ();
drwire add_88_21_n_951 ();
drwire add_88_21_n_953 ();
drwire add_88_21_n_955 ();
drwire add_88_21_n_957 ();
drwire add_88_21_n_979 ();
drwire add_88_21_n_980 ();
drwire add_88_21_n_982 ();
drwire add_88_21_n_985 ();
drwire add_88_21_n_987 ();
drwire add_88_21_n_989 ();
drwire add_88_21_n_991 ();
drwire add_88_21_n_992 ();
drwire add_88_21_n_996 ();
drwire add_88_21_n_997 ();
drwire add_88_21_n_999 ();
drwire add_88_69_n_1243 ();
drwire add_88_69_n_1259 ();
drwire add_88_69_n_1261 ();
drwire add_88_69_n_1262 ();
drwire add_88_69_n_1263 ();
drwire add_88_69_n_1265 ();
drwire add_88_69_n_1267 ();
drwire add_88_69_n_1268 ();
drwire add_88_69_n_1270 ();
drwire add_88_69_n_1271 ();
drwire add_88_69_n_1272 ();
drwire add_88_69_n_1274 ();
drwire add_88_69_n_1276 ();
drwire add_88_69_n_1277 ();
drwire add_88_69_n_1278 ();
drwire add_88_69_n_1280 ();
drwire add_88_69_n_1284 ();
drwire add_88_69_n_1288 ();
drwire add_88_69_n_1289 ();
drwire add_88_69_n_1290 ();
drwire add_88_69_n_1292 ();
drwire add_88_69_n_1293 ();
drwire add_88_69_n_1295 ();
drwire add_88_69_n_1297 ();
drwire add_88_69_n_1298 ();
drwire add_88_69_n_1300 ();
drwire add_88_69_n_1302 ();
drwire add_88_69_n_1303 ();
drwire add_88_69_n_1304 ();
drwire add_88_69_n_1308 ();
drwire add_88_69_n_1309 ();
drwire add_88_69_n_1311 ();
drwire add_88_69_n_1313 ();
drwire add_88_69_n_1315 ();
drwire add_88_69_n_1316 ();
drwire add_88_69_n_1318 ();
drwire add_88_69_n_1321 ();
drwire add_88_69_n_1322 ();
drwire add_88_69_n_1323 ();
drwire add_88_69_n_1327 ();
drwire add_88_69_n_1328 ();
drwire add_88_69_n_1329 ();
drwire add_88_69_n_1330 ();
drwire add_88_69_n_1331 ();
drwire add_88_69_n_1334 ();
drwire add_88_69_n_1337 ();
drwire add_88_69_n_1341 ();
drwire add_88_69_n_1342 ();
drwire add_88_69_n_1343 ();
drwire add_88_69_n_1344 ();
drwire add_88_69_n_1345 ();
drwire add_88_69_n_1347 ();
drwire add_88_69_n_1355 ();
drwire add_88_69_n_1356 ();
drwire add_88_69_n_1358 ();
drwire add_88_69_n_1359 ();
drwire add_88_69_n_1360 ();
drwire add_88_69_n_1363 ();
drwire add_88_69_n_1364 ();
drwire add_88_69_n_1366 ();
drwire add_88_69_n_1367 ();
drwire add_88_69_n_1368 ();
drwire add_88_69_n_1369 ();
drwire add_88_69_n_1370 ();
drwire add_88_69_n_1371 ();
drwire add_88_69_n_1372 ();
drwire add_88_69_n_1373 ();
drwire add_88_69_n_1376 ();
drwire add_88_69_n_1377 ();
drwire add_88_69_n_1378 ();
drwire add_88_69_n_1380 ();
drwire add_88_69_n_1381 ();
drwire add_88_69_n_1382 ();
drwire add_88_69_n_1385 ();
drwire add_88_69_n_1389 ();
drwire add_88_69_n_1395 ();
drwire add_88_69_n_1397 ();
drwire add_88_69_n_1398 ();
drwire add_88_69_n_1400 ();
drwire add_88_69_n_1404 ();
drwire add_88_69_n_1405 ();
drwire add_88_69_n_1406 ();
drwire add_88_69_n_1407 ();
drwire add_88_69_n_1408 ();
drwire add_88_69_n_1409 ();
drwire add_88_69_n_1412 ();
drwire add_88_69_n_1414 ();
drwire add_88_69_n_1417 ();
drwire add_88_69_n_1419 ();
drwire add_88_69_n_1422 ();
drwire add_88_69_n_1424 ();
drwire add_88_69_n_1425 ();
drwire add_88_69_n_1431 ();
drwire add_88_69_n_1437 ();
drwire add_88_69_n_1438 ();
drwire add_88_69_n_1439 ();
drwire add_88_69_n_1441 ();
drwire add_88_69_n_1443 ();
drwire add_88_69_n_1444 ();
drwire add_88_69_n_1445 ();
drwire add_88_69_n_1447 ();
drwire add_88_69_n_1449 ();
drwire add_88_69_n_1452 ();
drwire add_88_69_n_1453 ();
drwire add_88_69_n_1454 ();
drwire add_88_69_n_1456 ();
drwire add_88_69_n_1458 ();
drwire add_88_69_n_1464 ();
drwire add_88_69_n_1465 ();
drwire add_88_69_n_1466 ();
drwire add_88_69_n_1469 ();
drwire add_88_69_n_1470 ();
drwire add_88_69_n_1471 ();
drwire add_88_69_n_1472 ();
drwire add_88_69_n_1473 ();
drwire add_88_69_n_1474 ();
drwire add_88_69_n_1475 ();
drwire add_88_69_n_1476 ();
drwire add_88_69_n_1477 ();
drwire add_88_69_n_1478 ();
drwire add_88_69_n_1479 ();
drwire add_88_69_n_1481 ();
drwire add_88_69_n_1490 ();
drwire add_88_69_n_1491 ();
drwire add_88_69_n_1492 ();
drwire add_88_69_n_1496 ();
drwire add_88_69_n_1499 ();
drwire add_88_69_n_1500 ();
drwire add_88_69_n_1501 ();
drwire add_88_69_n_1502 ();
drwire add_88_69_n_1504 ();
drwire add_88_69_n_1505 ();
drwire add_88_69_n_1506 ();
drwire add_88_69_n_1508 ();
drwire add_88_69_n_1510 ();
drwire add_88_69_n_1513 ();
drwire add_88_69_n_1514 ();
drwire add_88_69_n_1515 ();
drwire add_88_69_n_1516 ();
drwire add_88_69_n_1518 ();
drwire add_88_69_n_1519 ();
drwire add_88_69_n_1520 ();
drwire add_88_69_n_1522 ();
drwire add_88_69_n_1523 ();
drwire add_88_69_n_1524 ();
drwire add_88_69_n_1525 ();
drwire add_88_69_n_1527 ();
drwire add_88_69_n_1528 ();
drwire add_88_69_n_1529 ();
drwire add_88_69_n_1530 ();
drwire add_88_69_n_1531 ();
drwire add_88_69_n_1532 ();
drwire add_88_69_n_1535 ();
drwire add_88_69_n_1536 ();
drwire add_88_69_n_1538 ();
drwire add_88_69_n_1543 ();
drwire add_88_69_n_1545 ();
drwire add_88_69_n_1547 ();
drwire add_88_69_n_1548 ();
drwire add_88_69_n_1551 ();
drwire add_88_69_n_1554 ();
drwire add_88_69_n_1556 ();
drwire add_88_69_n_1557 ();
drwire add_88_69_n_1601 ();
drwire add_88_69_n_1605 ();
drwire add_88_69_n_1606 ();
drwire add_88_69_n_1608 ();
drwire add_88_69_n_1612 ();
drwire add_88_69_n_1614 ();
drwire add_88_69_n_1631 ();
drwire add_88_69_n_1632 ();
drwire add_88_69_n_1633 ();
drwire add_88_69_n_1634 ();
drwire add_88_69_n_1635 ();
drwire add_88_69_n_1636 ();
drwire add_88_69_n_1638 ();
drwire add_88_69_n_1642 ();
drwire add_88_69_n_1643 ();
drwire add_88_69_n_1644 ();
drwire add_88_69_n_1645 ();
drwire add_88_69_n_1646 ();
drwire add_88_69_n_1647 ();
drwire add_88_69_n_1648 ();
drwire add_88_69_n_1649 ();
drwire add_88_69_n_1650 ();
drwire add_88_69_n_1653 ();
drwire add_88_69_n_1654 ();
drwire add_88_69_n_1655 ();
drwire add_88_69_n_1656 ();
drwire add_88_69_n_1659 ();
drwire add_88_69_n_1660 ();
drwire add_88_69_n_1662 ();
drwire add_88_69_n_1663 ();
drwire add_88_69_n_1668 ();
drwire add_88_69_n_1669 ();
drwire add_88_69_n_1670 ();
drwire add_88_69_n_1671 ();
drwire add_88_69_n_1672 ();
drwire add_88_69_n_1673 ();
drwire add_88_69_n_1674 ();
drwire add_88_69_n_1675 ();
drwire add_88_69_n_1676 ();
drwire add_88_69_n_1679 ();
drwire add_88_69_n_1680 ();
drwire add_88_69_n_1697 ();
drwire add_88_69_n_1698 ();
drwire add_88_69_n_1699 ();
drwire add_88_69_n_1700 ();
drwire add_88_69_n_1701 ();
drwire add_88_69_n_1702 ();
drwire add_88_69_n_1703 ();
drwire add_88_69_n_1704 ();
drwire add_88_69_n_1705 ();
drwire add_88_69_n_1706 ();
drwire add_88_69_n_1708 ();
drwire add_88_69_n_1709 ();
drwire add_88_69_n_1710 ();
drwire add_88_69_n_1711 ();
drwire add_88_69_n_1712 ();
drwire add_88_69_n_1714 ();
drwire add_88_69_n_1715 ();
drwire add_88_69_n_1716 ();
drwire add_88_69_n_1717 ();
drwire add_88_69_n_1718 ();
drwire add_88_69_n_1719 ();
drwire add_88_69_n_1720 ();
drwire add_88_69_n_1721 ();
drwire add_88_69_n_1722 ();
drwire add_88_69_n_1723 ();
drwire add_88_69_n_1725 ();
drwire add_88_69_n_1727 ();
drwire add_88_69_n_1728 ();
drwire add_88_69_n_1729 ();
drwire add_88_69_n_1730 ();
drwire add_88_69_n_1731 ();
drwire add_88_69_n_1732 ();
drwire add_88_69_n_1734 ();
drwire add_88_69_n_1735 ();
drwire add_88_69_n_1736 ();
drwire add_88_69_n_1737 ();
drwire add_88_69_n_1739 ();
drwire add_88_69_n_1740 ();
drwire add_88_69_n_1741 ();
drwire add_88_69_n_1743 ();
drwire add_88_69_n_1745 ();
drwire add_88_69_n_1746 ();
drwire add_88_69_n_1749 ();
drwire add_88_69_n_1752 ();
drwire add_88_69_n_1755 ();
drwire add_88_82_n_1889 ();
drwire add_88_82_n_1893 ();
drwire add_88_82_n_1896 ();
drwire add_88_82_n_1899 ();
drwire add_88_82_n_1900 ();
drwire add_88_82_n_1903 ();
drwire add_88_82_n_1905 ();
drwire add_88_82_n_1906 ();
drwire add_88_82_n_1910 ();
drwire add_88_82_n_1911 ();
drwire add_88_82_n_1913 ();
drwire add_88_82_n_1917 ();
drwire add_88_82_n_1918 ();
drwire add_88_82_n_1920 ();
drwire add_88_82_n_1921 ();
drwire add_88_82_n_1925 ();
drwire add_88_82_n_1926 ();
drwire add_88_82_n_1928 ();
drwire add_88_82_n_1930 ();
drwire add_88_82_n_1932 ();
drwire add_88_82_n_1936 ();
drwire add_88_82_n_1938 ();
drwire add_88_82_n_1939 ();
drwire add_88_82_n_1940 ();
drwire add_88_82_n_1941 ();
drwire add_88_82_n_1945 ();
drwire add_88_82_n_1947 ();
drwire add_88_82_n_1949 ();
drwire add_88_82_n_1950 ();
drwire add_88_82_n_1952 ();
drwire add_88_82_n_1958 ();
drwire add_88_82_n_1959 ();
drwire add_88_82_n_1960 ();
drwire add_88_82_n_1961 ();
drwire add_88_82_n_1965 ();
drwire add_88_82_n_1967 ();
drwire add_88_82_n_1968 ();
drwire add_88_82_n_1969 ();
drwire add_88_82_n_1971 ();
drwire add_88_82_n_1973 ();
drwire add_88_82_n_1974 ();
drwire add_88_82_n_1975 ();
drwire add_88_82_n_1977 ();
drwire add_88_82_n_1978 ();
drwire add_88_82_n_1981 ();
drwire add_88_82_n_1982 ();
drwire add_88_82_n_1985 ();
drwire add_88_82_n_1987 ();
drwire add_88_82_n_1988 ();
drwire add_88_82_n_1989 ();
drwire add_88_82_n_1991 ();
drwire add_88_82_n_1993 ();
drwire add_88_82_n_1994 ();
drwire add_88_82_n_1996 ();
drwire add_88_82_n_1997 ();
drwire add_88_82_n_1999 ();
drwire add_88_82_n_2001 ();
drwire add_88_82_n_2003 ();
drwire add_88_82_n_2004 ();
drwire add_88_82_n_2005 ();
drwire add_88_82_n_2006 ();
drwire add_88_82_n_2007 ();
drwire add_88_82_n_2008 ();
drwire add_88_82_n_2010 ();
drwire add_88_82_n_2011 ();
drwire add_88_82_n_2013 ();
drwire add_88_82_n_2014 ();
drwire add_88_82_n_2015 ();
drwire add_88_82_n_2016 ();
drwire add_88_82_n_2018 ();
drwire add_88_82_n_2020 ();
drwire add_88_82_n_2023 ();
drwire add_88_82_n_2024 ();
drwire add_88_82_n_2025 ();
drwire add_88_82_n_2026 ();
drwire add_88_82_n_2027 ();
drwire add_88_82_n_2028 ();
drwire add_88_82_n_2029 ();
drwire add_88_82_n_2030 ();
drwire add_88_82_n_2034 ();
drwire add_88_82_n_2035 ();
drwire add_88_82_n_2037 ();
drwire add_88_82_n_2038 ();
drwire add_88_82_n_2039 ();
drwire add_88_82_n_2040 ();
drwire add_88_82_n_2041 ();
drwire add_88_82_n_2042 ();
drwire add_88_82_n_2044 ();
drwire add_88_82_n_2045 ();
drwire add_88_82_n_2048 ();
drwire add_88_82_n_2050 ();
drwire add_88_82_n_2051 ();
drwire add_88_82_n_2052 ();
drwire add_88_82_n_2053 ();
drwire add_88_82_n_2054 ();
drwire add_88_82_n_2055 ();
drwire add_88_82_n_2056 ();
drwire add_88_82_n_2057 ();
drwire add_88_82_n_2058 ();
drwire add_88_82_n_2059 ();
drwire add_88_82_n_2060 ();
drwire add_88_82_n_2061 ();
drwire add_88_82_n_2062 ();
drwire add_88_82_n_2063 ();
drwire add_88_82_n_2064 ();
drwire add_88_82_n_2065 ();
drwire add_88_82_n_2067 ();
drwire add_88_82_n_2069 ();
drwire add_88_82_n_2074 ();
drwire add_88_82_n_2076 ();
drwire add_88_82_n_2078 ();
drwire add_88_82_n_2079 ();
drwire add_88_82_n_2081 ();
drwire add_88_82_n_2082 ();
drwire add_88_82_n_2084 ();
drwire add_88_82_n_2086 ();
drwire add_88_82_n_2088 ();
drwire add_88_82_n_2091 ();
drwire add_88_82_n_2093 ();
drwire add_88_82_n_2096 ();
drwire add_88_82_n_2099 ();
drwire add_88_82_n_2101 ();
drwire add_88_82_n_2103 ();
drwire add_88_82_n_2105 ();
drwire add_88_82_n_2107 ();
drwire add_88_82_n_2109 ();
drwire add_88_82_n_2110 ();
drwire add_88_82_n_2111 ();
drwire add_88_82_n_2116 ();
drwire add_88_82_n_2117 ();
drwire add_88_82_n_2118 ();
drwire add_88_82_n_2120 ();
drwire add_88_82_n_2121 ();
drwire add_88_82_n_2122 ();
drwire add_88_82_n_2123 ();
drwire add_88_82_n_2124 ();
drwire add_88_82_n_2125 ();
drwire add_88_82_n_2126 ();
drwire add_88_82_n_2127 ();
drwire add_88_82_n_2128 ();
drwire add_88_82_n_2129 ();
drwire add_88_82_n_2130 ();
drwire add_88_82_n_2131 ();
drwire add_88_82_n_2132 ();
drwire add_88_82_n_2133 ();
drwire add_88_82_n_2134 ();
drwire add_88_82_n_2135 ();
drwire add_88_82_n_2136 ();
drwire add_88_82_n_2137 ();
drwire add_88_82_n_2138 ();
drwire add_88_82_n_2139 ();
drwire add_88_82_n_2141 ();
drwire add_88_82_n_2142 ();
drwire add_88_82_n_2143 ();
drwire add_88_82_n_2144 ();
drwire add_88_82_n_2145 ();
drwire add_88_82_n_2146 ();
drwire add_88_82_n_2147 ();
drwire add_88_82_n_2148 ();
drwire add_88_82_n_2149 ();
drwire add_88_82_n_2152 ();
drwire add_88_82_n_2153 ();
drwire add_88_82_n_2154 ();
drwire add_88_82_n_2155 ();
drwire add_88_82_n_2156 ();
drwire add_88_82_n_2157 ();
drwire add_88_82_n_2158 ();
drwire add_88_82_n_2159 ();
drwire add_88_82_n_2160 ();
drwire add_88_82_n_2161 ();
drwire add_88_82_n_2162 ();
drwire add_88_82_n_2163 ();
drwire add_88_82_n_2164 ();
drwire add_88_82_n_2165 ();
drwire add_88_82_n_2166 ();
drwire add_88_82_n_2167 ();
drwire add_88_82_n_2168 ();
drwire add_88_82_n_2169 ();
drwire add_88_82_n_2170 ();
drwire add_88_82_n_2171 ();
drwire add_88_82_n_2172 ();
drwire add_88_82_n_2173 ();
drwire add_88_82_n_2174 ();
drwire add_88_82_n_2176 ();
drwire add_88_82_n_2177 ();
drwire add_88_82_n_2178 ();
drwire add_88_82_n_2179 ();
drwire add_88_82_n_2180 ();
drwire add_88_82_n_2181 ();
drwire add_88_82_n_2182 ();
drwire add_88_82_n_2185 ();
drwire add_88_82_n_2188 ();
drwire add_88_82_n_2189 ();
drwire add_88_82_n_2190 ();
drwire add_88_82_n_2193 ();
drwire add_88_82_n_2196 ();
drwire add_88_82_n_2199 ();
drwire add_88_82_n_2202 ();
drwire add_88_82_n_2208 ();
drwire add_88_82_n_2231 ();
drwire add_88_82_n_2235 ();
drwire add_88_82_n_2236 ();
drwire add_88_82_n_2237 ();
drwire add_88_82_n_2238 ();
drwire add_88_82_n_2239 ();
drwire add_88_82_n_2241 ();
drwire add_88_82_n_2242 ();
drwire add_88_82_n_2243 ();
drwire add_88_82_n_2244 ();
drwire add_88_82_n_2245 ();
drwire add_88_82_n_2246 ();
drwire add_88_82_n_2247 ();
drwire add_88_82_n_2248 ();
drwire add_88_82_n_2249 ();
drwire add_88_82_n_2250 ();
drwire add_88_82_n_2251 ();
drwire add_88_82_n_2252 ();
drwire add_88_82_n_2253 ();
drwire add_88_82_n_2254 ();
drwire add_88_82_n_2255 ();
drwire add_88_82_n_2256 ();
drwire add_88_82_n_2257 ();
drwire add_88_82_n_2258 ();
drwire add_88_82_n_2259 ();
drwire add_88_82_n_2260 ();
drwire add_88_82_n_2261 ();
drwire add_88_82_n_2262 ();
drwire add_88_82_n_2263 ();
drwire add_88_82_n_2264 ();
drwire add_88_82_n_2265 ();
drwire add_88_82_n_2266 ();
drwire add_88_82_n_2267 ();
drwire add_88_82_n_2268 ();
drwire add_88_82_n_2269 ();
drwire add_88_82_n_2270 ();
drwire add_88_82_n_2271 ();
drwire add_88_82_n_2274 ();
drwire add_88_82_n_2277 ();
drwire add_88_82_n_2280 ();
drwire add_88_82_n_2283 ();
drwire add_88_82_n_2286 ();
drwire add_88_82_n_2287 ();
drwire add_88_82_n_2288 ();
drwire add_88_82_n_2289 ();
drwire add_88_82_n_2292 ();
drwire add_88_82_n_2293 ();
drwire add_88_82_n_2371 ();
drwire add_88_82_n_2372 ();
drwire counter_10_ ();
drwire counter_1_ ();
drwire counter_2_ ();
drwire counter_3_ ();
drwire counter_4_ ();
drwire counter_5_ ();
drwire counter_6_ ();
drwire counter_7_ ();
drwire counter_8_ ();
drwire counter_9_ ();
drwire inc_add_77_23_n_411 ();
drwire inc_add_77_23_n_412 ();
drwire inc_add_77_23_n_413 ();
drwire inc_add_77_23_n_421 ();
drwire inc_add_77_23_n_422 ();
drwire inc_add_77_23_n_424 ();
drwire inc_add_77_23_n_426 ();
drwire inc_add_77_23_n_427 ();
drwire inc_add_77_23_n_428 ();
drwire inc_add_77_23_n_430 ();
drwire inc_add_77_23_n_431 ();
drwire inc_add_77_23_n_432 ();
drwire inc_add_77_23_n_433 ();
drwire inc_add_77_23_n_435 ();
drwire inc_add_77_23_n_439 ();
drwire inc_add_77_23_n_440 ();
drwire inc_add_77_23_n_441 ();
drwire inc_add_77_23_n_442 ();
drwire inc_add_77_23_n_443 ();
drwire inc_add_77_23_n_444 ();
drwire inc_add_77_23_n_445 ();
drwire inc_add_77_23_n_446 ();
drwire inc_add_77_23_n_448 ();
drwire inc_add_77_23_n_451 ();
drwire inc_add_77_23_n_453 ();
drwire inc_add_77_23_n_454 ();
drwire inc_add_77_23_n_455 ();
drwire inc_add_77_23_n_458 ();
drwire inc_add_77_23_n_460 ();
drwire inc_add_77_23_n_462 ();
drwire inc_add_77_23_n_463 ();
drwire inc_add_77_23_n_464 ();
drwire inc_add_77_23_n_465 ();
drwire inc_add_77_23_n_469 ();
drwire inc_add_77_23_n_470 ();
drwire inc_add_77_23_n_476 ();
drwire inc_add_77_23_n_478 ();
drwire inc_add_77_23_n_482 ();
drwire inc_add_77_23_n_483 ();
drwire inc_add_77_23_n_484 ();
drwire inc_add_77_23_n_485 ();
drwire inc_add_77_23_n_486 ();
drwire inc_add_77_23_n_487 ();
drwire inc_add_77_23_n_489 ();
drwire inc_add_77_23_n_490 ();
drwire inc_add_77_23_n_491 ();
drwire inc_add_77_23_n_492 ();
drwire inc_add_77_23_n_493 ();
drwire inc_add_77_23_n_494 ();
drwire inc_add_77_23_n_495 ();
drwire inc_add_77_23_n_496 ();
drwire inc_add_77_23_n_498 ();
drwire inc_add_77_23_n_501 ();
drwire inc_add_77_23_n_502 ();
drwire inc_add_77_23_n_506 ();
drwire inc_add_77_23_n_508 ();
drwire inc_add_77_23_n_510 ();
drwire inc_add_77_23_n_512 ();
drwire inc_add_77_23_n_515 ();
drwire inc_add_77_23_n_517 ();
drwire inc_add_77_23_n_520 ();
drwire inc_add_77_23_n_522 ();
drwire inc_add_77_23_n_523 ();
drwire inc_add_77_23_n_524 ();
drwire inc_add_77_23_n_525 ();
drwire inc_add_77_23_n_526 ();
drwire inc_add_77_23_n_527 ();
drwire inc_add_77_23_n_528 ();
drwire inc_add_77_23_n_530 ();
drwire inc_add_77_23_n_532 ();
drwire inc_add_77_23_n_540 ();
drwire inc_add_77_23_n_541 ();
drwire inc_add_77_23_n_542 ();
drwire inc_add_77_23_n_543 ();
drwire inc_add_77_23_n_544 ();
drwire inc_add_77_23_n_545 ();
drwire inc_add_77_23_n_546 ();
drwire inc_add_77_23_n_547 ();
drwire inc_add_77_23_n_549 ();
drwire inc_add_77_23_n_551 ();
drwire inc_add_77_23_n_553 ();
drwire inc_add_77_23_n_562 ();
drwire inc_add_77_23_n_566 ();
drwire inc_add_77_23_n_569 ();
drwire inc_add_77_23_n_572 ();
drwire inc_add_77_23_n_581 ();
drwire inc_add_77_23_n_585 ();
drwire inc_add_77_23_n_591 ();
drwire inc_add_77_23_n_593 ();
drwire key_r_0_ ();
drwire key_r_100_ ();
drwire key_r_101_ ();
drwire key_r_102_ ();
drwire key_r_103_ ();
drwire key_r_104_ ();
drwire key_r_105_ ();
drwire key_r_106_ ();
drwire key_r_107_ ();
drwire key_r_108_ ();
drwire key_r_109_ ();
drwire key_r_10_ ();
drwire key_r_110_ ();
drwire key_r_111_ ();
drwire key_r_112_ ();
drwire key_r_113_ ();
drwire key_r_114_ ();
drwire key_r_115_ ();
drwire key_r_116_ ();
drwire key_r_117_ ();
drwire key_r_118_ ();
drwire key_r_119_ ();
drwire key_r_11_ ();
drwire key_r_120_ ();
drwire key_r_121_ ();
drwire key_r_122_ ();
drwire key_r_123_ ();
drwire key_r_124_ ();
drwire key_r_125_ ();
drwire key_r_126_ ();
drwire key_r_127_ ();
drwire key_r_12_ ();
drwire key_r_13_ ();
drwire key_r_14_ ();
drwire key_r_15_ ();
drwire key_r_16_ ();
drwire key_r_17_ ();
drwire key_r_18_ ();
drwire key_r_19_ ();
drwire key_r_1_ ();
drwire key_r_20_ ();
drwire key_r_21_ ();
drwire key_r_22_ ();
drwire key_r_23_ ();
drwire key_r_24_ ();
drwire key_r_25_ ();
drwire key_r_26_ ();
drwire key_r_27_ ();
drwire key_r_28_ ();
drwire key_r_29_ ();
drwire key_r_2_ ();
drwire key_r_30_ ();
drwire key_r_31_ ();
drwire key_r_32_ ();
drwire key_r_33_ ();
drwire key_r_34_ ();
drwire key_r_35_ ();
drwire key_r_36_ ();
drwire key_r_37_ ();
drwire key_r_38_ ();
drwire key_r_39_ ();
drwire key_r_3_ ();
drwire key_r_40_ ();
drwire key_r_41_ ();
drwire key_r_42_ ();
drwire key_r_43_ ();
drwire key_r_44_ ();
drwire key_r_45_ ();
drwire key_r_46_ ();
drwire key_r_47_ ();
drwire key_r_48_ ();
drwire key_r_49_ ();
drwire key_r_4_ ();
drwire key_r_50_ ();
drwire key_r_51_ ();
drwire key_r_52_ ();
drwire key_r_53_ ();
drwire key_r_54_ ();
drwire key_r_55_ ();
drwire key_r_56_ ();
drwire key_r_57_ ();
drwire key_r_58_ ();
drwire key_r_59_ ();
drwire key_r_5_ ();
drwire key_r_60_ ();
drwire key_r_61_ ();
drwire key_r_62_ ();
drwire key_r_63_ ();
drwire key_r_64_ ();
drwire key_r_65_ ();
drwire key_r_66_ ();
drwire key_r_67_ ();
drwire key_r_68_ ();
drwire key_r_69_ ();
drwire key_r_6_ ();
drwire key_r_70_ ();
drwire key_r_71_ ();
drwire key_r_72_ ();
drwire key_r_73_ ();
drwire key_r_74_ ();
drwire key_r_75_ ();
drwire key_r_76_ ();
drwire key_r_77_ ();
drwire key_r_78_ ();
drwire key_r_79_ ();
drwire key_r_7_ ();
drwire key_r_80_ ();
drwire key_r_81_ ();
drwire key_r_82_ ();
drwire key_r_83_ ();
drwire key_r_84_ ();
drwire key_r_85_ ();
drwire key_r_86_ ();
drwire key_r_87_ ();
drwire key_r_88_ ();
drwire key_r_89_ ();
drwire key_r_8_ ();
drwire key_r_90_ ();
drwire key_r_91_ ();
drwire key_r_92_ ();
drwire key_r_93_ ();
drwire key_r_94_ ();
drwire key_r_95_ ();
drwire key_r_96_ ();
drwire key_r_97_ ();
drwire key_r_98_ ();
drwire key_r_99_ ();
drwire key_r_9_ ();
drwire n_0 ();
drwire n_1 ();
drwire n_100 ();
drwire n_101 ();
drwire n_11 ();
drwire n_117 ();
drwire n_12 ();
drwire n_1216 ();
drwire n_1217 ();
drwire n_1224 ();
drwire n_1235 ();
drwire n_1239 ();
drwire n_1240 ();
drwire n_1241 ();
drwire n_1243 ();
drwire n_1244 ();
drwire n_1245 ();
drwire n_1246 ();
drwire n_125 ();
drwire n_128 ();
drwire n_1280 ();
drwire n_1281 ();
drwire n_1282 ();
drwire n_1283 ();
drwire n_1284 ();
drwire n_1285 ();
drwire n_1286 ();
drwire n_1287 ();
drwire n_1288 ();
drwire n_1289 ();
drwire n_129 ();
drwire n_1290 ();
drwire n_1291 ();
drwire n_1292 ();
drwire n_1293 ();
drwire n_1294 ();
drwire n_1295 ();
drwire n_1296 ();
drwire n_1297 ();
drwire n_1298 ();
drwire n_13 ();
drwire n_1301 ();
drwire n_1302 ();
drwire n_1303 ();
drwire n_1304 ();
drwire n_1305 ();
drwire n_1306 ();
drwire n_1307 ();
drwire n_1308 ();
drwire n_131 ();
drwire n_1312 ();
drwire n_1313 ();
drwire n_1314 ();
drwire n_1315 ();
drwire n_1316 ();
drwire n_132 ();
drwire n_1322 ();
drwire n_1323 ();
drwire n_133 ();
drwire n_1330 ();
drwire n_134 ();
drwire n_1345 ();
drwire n_1346 ();
drwire n_1347 ();
drwire n_1348 ();
drwire n_135 ();
drwire n_1359 ();
drwire n_136 ();
drwire n_1360 ();
drwire n_1361 ();
drwire n_1362 ();
drwire n_137 ();
drwire n_1379 ();
drwire n_138 ();
drwire n_1386 ();
drwire n_1387 ();
drwire n_1388 ();
drwire n_1389 ();
drwire n_139 ();
drwire n_1393 ();
drwire n_14 ();
drwire n_140 ();
drwire n_1400 ();
drwire n_1407 ();
drwire n_141 ();
drwire n_1414 ();
drwire n_142 ();
drwire n_1421 ();
drwire n_1428 ();
drwire n_143 ();
drwire n_144 ();
drwire n_1442 ();
drwire n_1443 ();
drwire n_1444 ();
drwire n_1445 ();
drwire n_1446 ();
drwire n_1447 ();
drwire n_1449 ();
drwire n_145 ();
drwire n_1450 ();
drwire n_1451 ();
drwire n_1452 ();
drwire n_1453 ();
drwire n_1459 ();
drwire n_146 ();
drwire n_1463 ();
drwire n_1464 ();
drwire n_1465 ();
drwire n_1469 ();
drwire n_147 ();
drwire n_1470 ();
drwire n_1471 ();
drwire n_1472 ();
drwire n_1473 ();
drwire n_1475 ();
drwire n_1476 ();
drwire n_1477 ();
drwire n_1478 ();
drwire n_1479 ();
drwire n_148 ();
drwire n_1481 ();
drwire n_1483 ();
drwire n_1484 ();
drwire n_1487 ();
drwire n_1488 ();
drwire n_1489 ();
drwire n_149 ();
drwire n_1490 ();
drwire n_1494 ();
drwire n_1495 ();
drwire n_1496 ();
drwire n_1497 ();
drwire n_1498 ();
drwire n_15 ();
drwire n_150 ();
drwire n_1500 ();
drwire n_1501 ();
drwire n_1502 ();
drwire n_1503 ();
drwire n_1504 ();
drwire n_1507 ();
drwire n_1508 ();
drwire n_1509 ();
drwire n_151 ();
drwire n_1510 ();
drwire n_1511 ();
drwire n_1512 ();
drwire n_1513 ();
drwire n_1514 ();
drwire n_1515 ();
drwire n_1516 ();
drwire n_1517 ();
drwire n_152 ();
drwire n_1526 ();
drwire n_1527 ();
drwire n_1528 ();
drwire n_153 ();
drwire n_1538 ();
drwire n_1539 ();
drwire n_154 ();
drwire n_1540 ();
drwire n_1541 ();
drwire n_1544 ();
drwire n_1548 ();
drwire n_1550 ();
drwire n_1551 ();
drwire n_1552 ();
drwire n_1553 ();
drwire n_1554 ();
drwire n_1555 ();
drwire n_1556 ();
drwire n_1557 ();
drwire n_156 ();
drwire n_1561 ();
drwire n_1563 ();
drwire n_1564 ();
drwire n_157 ();
drwire n_1572 ();
drwire n_1573 ();
drwire n_1574 ();
drwire n_1578 ();
drwire n_1579 ();
drwire n_158 ();
drwire n_1580 ();
drwire n_1584 ();
drwire n_1585 ();
drwire n_1586 ();
drwire n_1587 ();
drwire n_1588 ();
drwire n_1589 ();
drwire n_159 ();
drwire n_1590 ();
drwire n_1591 ();
drwire n_1592 ();
drwire n_1593 ();
drwire n_1594 ();
drwire n_1595 ();
drwire n_1596 ();
drwire n_1597 ();
drwire n_1598 ();
drwire n_16 ();
drwire n_160 ();
drwire n_1605 ();
drwire n_1606 ();
drwire n_1607 ();
drwire n_1608 ();
drwire n_161 ();
drwire n_1619 ();
drwire n_162 ();
drwire n_1620 ();
drwire n_1621 ();
drwire n_1622 ();
drwire n_1623 ();
drwire n_1624 ();
drwire n_1625 ();
drwire n_1626 ();
drwire n_1627 ();
drwire n_1628 ();
drwire n_1629 ();
drwire n_163 ();
drwire n_1630 ();
drwire n_1631 ();
drwire n_1633 ();
drwire n_1635 ();
drwire n_1636 ();
drwire n_1637 ();
drwire n_1638 ();
drwire n_1639 ();
drwire n_164 ();
drwire n_1640 ();
drwire n_1641 ();
drwire n_1642 ();
drwire n_1643 ();
drwire n_1644 ();
drwire n_1645 ();
drwire n_1646 ();
drwire n_1647 ();
drwire n_165 ();
drwire n_1651 ();
drwire n_1652 ();
drwire n_1653 ();
drwire n_1654 ();
drwire n_1655 ();
drwire n_1656 ();
drwire n_1658 ();
drwire n_166 ();
drwire n_1660 ();
drwire n_1661 ();
drwire n_1662 ();
drwire n_1663 ();
drwire n_1664 ();
drwire n_1665 ();
drwire n_1666 ();
drwire n_1667 ();
drwire n_1668 ();
drwire n_167 ();
drwire n_1670 ();
drwire n_1671 ();
drwire n_1672 ();
drwire n_1673 ();
drwire n_1674 ();
drwire n_1676 ();
drwire n_1677 ();
drwire n_1678 ();
drwire n_168 ();
drwire n_1681 ();
drwire n_1682 ();
drwire n_1683 ();
drwire n_1684 ();
drwire n_1685 ();
drwire n_1686 ();
drwire n_1687 ();
drwire n_1688 ();
drwire n_1689 ();
drwire n_169 ();
drwire n_1690 ();
drwire n_1691 ();
drwire n_1698 ();
drwire n_1699 ();
drwire n_17 ();
drwire n_170 ();
drwire n_1700 ();
drwire n_1701 ();
drwire n_1702 ();
drwire n_1703 ();
drwire n_1704 ();
drwire n_1705 ();
drwire n_1706 ();
drwire n_1707 ();
drwire n_1709 ();
drwire n_171 ();
drwire n_1710 ();
drwire n_1711 ();
drwire n_1712 ();
drwire n_1713 ();
drwire n_1714 ();
drwire n_1718 ();
drwire n_1719 ();
drwire n_172 ();
drwire n_1721 ();
drwire n_1722 ();
drwire n_1723 ();
drwire n_1724 ();
drwire n_1725 ();
drwire n_1726 ();
drwire n_1727 ();
drwire n_1728 ();
drwire n_1729 ();
drwire n_173 ();
drwire n_1730 ();
drwire n_1731 ();
drwire n_1732 ();
drwire n_1733 ();
drwire n_1737 ();
drwire n_174 ();
drwire n_1740 ();
drwire n_1741 ();
drwire n_1742 ();
drwire n_1745 ();
drwire n_1746 ();
drwire n_1747 ();
drwire n_1748 ();
drwire n_1749 ();
drwire n_175 ();
drwire n_1750 ();
drwire n_1751 ();
drwire n_1752 ();
drwire n_1753 ();
drwire n_1754 ();
drwire n_1755 ();
drwire n_1756 ();
drwire n_1757 ();
drwire n_1758 ();
drwire n_1762 ();
drwire n_1764 ();
drwire n_1765 ();
drwire n_1766 ();
drwire n_1769 ();
drwire n_1771 ();
drwire n_1772 ();
drwire n_1773 ();
drwire n_1774 ();
drwire n_1775 ();
drwire n_1776 ();
drwire n_1779 ();
drwire n_178 ();
drwire n_1782 ();
drwire n_1785 ();
drwire n_1789 ();
drwire n_179 ();
drwire n_1791 ();
drwire n_1792 ();
drwire n_1793 ();
drwire n_1794 ();
drwire n_1795 ();
drwire n_1796 ();
drwire n_1797 ();
drwire n_18 ();
drwire n_180 ();
drwire n_1800 ();
drwire n_1803 ();
drwire n_1804 ();
drwire n_1805 ();
drwire n_1806 ();
drwire n_1807 ();
drwire n_1808 ();
drwire n_181 ();
drwire n_1810 ();
drwire n_1812 ();
drwire n_1813 ();
drwire n_1815 ();
drwire n_1816 ();
drwire n_1817 ();
drwire n_1818 ();
drwire n_1819 ();
drwire n_182 ();
drwire n_1820 ();
drwire n_1827 ();
drwire n_1841 ();
drwire n_1842 ();
drwire n_1843 ();
drwire n_1844 ();
drwire n_1845 ();
drwire n_1846 ();
drwire n_1848 ();
drwire n_1849 ();
drwire n_1850 ();
drwire n_1859 ();
drwire n_1860 ();
drwire n_1861 ();
drwire n_1862 ();
drwire n_1866 ();
drwire n_1867 ();
drwire n_1868 ();
drwire n_1869 ();
drwire n_187 ();
drwire n_1870 ();
drwire n_1881 ();
drwire n_1882 ();
drwire n_1884 ();
drwire n_1885 ();
drwire n_1886 ();
drwire n_1887 ();
drwire n_1888 ();
drwire n_1889 ();
drwire n_1890 ();
drwire n_1892 ();
drwire n_1894 ();
drwire n_1895 ();
drwire n_19 ();
drwire n_1904 ();
drwire n_1905 ();
drwire n_1906 ();
drwire n_191 ();
drwire n_1910 ();
drwire n_1914 ();
drwire n_1915 ();
drwire n_1916 ();
drwire n_1917 ();
drwire n_1918 ();
drwire n_1919 ();
drwire n_192 ();
drwire n_1921 ();
drwire n_1922 ();
drwire n_1924 ();
drwire n_1927 ();
drwire n_1928 ();
drwire n_1929 ();
drwire n_193 ();
drwire n_1930 ();
drwire n_1931 ();
drwire n_1935 ();
drwire n_1936 ();
drwire n_194 ();
drwire n_1941 ();
drwire n_1946 ();
drwire n_1948 ();
drwire n_1950 ();
drwire n_1952 ();
drwire n_1954 ();
drwire n_1955 ();
drwire n_1956 ();
drwire n_1959 ();
drwire n_196 ();
drwire n_1962 ();
drwire n_1963 ();
drwire n_1964 ();
drwire n_1966 ();
drwire n_1967 ();
drwire n_1968 ();
drwire n_1969 ();
drwire n_1970 ();
drwire n_1971 ();
drwire n_1977 ();
drwire n_198 ();
drwire n_1980 ();
drwire n_1983 ();
drwire n_1984 ();
drwire n_1985 ();
drwire n_1986 ();
drwire n_1987 ();
drwire n_1989 ();
drwire n_1990 ();
drwire n_1991 ();
drwire n_1996 ();
drwire n_1997 ();
drwire n_1998 ();
drwire n_20 ();
drwire n_200 ();
drwire n_2003 ();
drwire n_2004 ();
drwire n_2005 ();
drwire n_2007 ();
drwire n_2014 ();
drwire n_2017 ();
drwire n_2018 ();
drwire n_2019 ();
drwire n_202 ();
drwire n_2020 ();
drwire n_2025 ();
drwire n_2026 ();
drwire n_2027 ();
drwire n_2028 ();
drwire n_2029 ();
drwire n_2030 ();
drwire n_2031 ();
drwire n_2033 ();
drwire n_2034 ();
drwire n_2035 ();
drwire n_2036 ();
drwire n_2037 ();
drwire n_2038 ();
drwire n_2039 ();
drwire n_2041 ();
drwire n_2042 ();
drwire n_2043 ();
drwire n_2044 ();
drwire n_2045 ();
drwire n_2049 ();
drwire n_205 ();
drwire n_2054 ();
drwire n_2057 ();
drwire n_2058 ();
drwire n_206 ();
drwire n_2060 ();
drwire n_2062 ();
drwire n_2063 ();
drwire n_2064 ();
drwire n_2065 ();
drwire n_2066 ();
drwire n_2067 ();
drwire n_2068 ();
drwire n_2069 ();
drwire n_207 ();
drwire n_2070 ();
drwire n_2071 ();
drwire n_2072 ();
drwire n_2073 ();
drwire n_2074 ();
drwire n_2075 ();
drwire n_2076 ();
drwire n_2077 ();
drwire n_2078 ();
drwire n_2079 ();
drwire n_208 ();
drwire n_2080 ();
drwire n_2085 ();
drwire n_2089 ();
drwire n_2091 ();
drwire n_2092 ();
drwire n_2096 ();
drwire n_2099 ();
drwire n_21 ();
drwire n_2100 ();
drwire n_2101 ();
drwire n_2102 ();
drwire n_2103 ();
drwire n_2104 ();
drwire n_2105 ();
drwire n_2106 ();
drwire n_2107 ();
drwire n_2108 ();
drwire n_2109 ();
drwire n_211 ();
drwire n_2110 ();
drwire n_2111 ();
drwire n_2112 ();
drwire n_2113 ();
drwire n_2115 ();
drwire n_2116 ();
drwire n_2117 ();
drwire n_2118 ();
drwire n_2119 ();
drwire n_212 ();
drwire n_2120 ();
drwire n_2121 ();
drwire n_2122 ();
drwire n_2123 ();
drwire n_2124 ();
drwire n_2125 ();
drwire n_2126 ();
drwire n_213 ();
drwire n_2131 ();
drwire n_2133 ();
drwire n_2134 ();
drwire n_2135 ();
drwire n_2136 ();
drwire n_2137 ();
drwire n_2138 ();
drwire n_214 ();
drwire n_2140 ();
drwire n_2142 ();
drwire n_2144 ();
drwire n_2145 ();
drwire n_2147 ();
drwire n_2149 ();
drwire n_215 ();
drwire n_2151 ();
drwire n_2152 ();
drwire n_2154 ();
drwire n_2156 ();
drwire n_2158 ();
drwire n_2159 ();
drwire n_216 ();
drwire n_2161 ();
drwire n_2163 ();
drwire n_2165 ();
drwire n_2166 ();
drwire n_2168 ();
drwire n_217 ();
drwire n_2170 ();
drwire n_2172 ();
drwire n_2173 ();
drwire n_2175 ();
drwire n_2177 ();
drwire n_2179 ();
drwire n_218 ();
drwire n_2182 ();
drwire n_2184 ();
drwire n_2186 ();
drwire n_2187 ();
drwire n_2189 ();
drwire n_219 ();
drwire n_2191 ();
drwire n_2193 ();
drwire n_2194 ();
drwire n_2195 ();
drwire n_2196 ();
drwire n_2197 ();
drwire n_2198 ();
drwire n_2199 ();
drwire n_220 ();
drwire n_2200 ();
drwire n_2201 ();
drwire n_2202 ();
drwire n_2204 ();
drwire n_221 ();
drwire n_2211 ();
drwire n_2212 ();
drwire n_2213 ();
drwire n_2214 ();
drwire n_2215 ();
drwire n_2216 ();
drwire n_2217 ();
drwire n_2218 ();
drwire n_2219 ();
drwire n_222 ();
drwire n_2222 ();
drwire n_2223 ();
drwire n_2224 ();
drwire n_2225 ();
drwire n_2226 ();
drwire n_2227 ();
drwire n_2228 ();
drwire n_2229 ();
drwire n_223 ();
drwire n_2230 ();
drwire n_2231 ();
drwire n_2232 ();
drwire n_2233 ();
drwire n_2235 ();
drwire n_2236 ();
drwire n_2237 ();
drwire n_224 ();
drwire n_2246 ();
drwire n_2247 ();
drwire n_225 ();
drwire n_2250 ();
drwire n_2251 ();
drwire n_2254 ();
drwire n_2255 ();
drwire n_2256 ();
drwire n_226 ();
drwire n_2261 ();
drwire n_2262 ();
drwire n_2269 ();
drwire n_227 ();
drwire n_2270 ();
drwire n_2271 ();
drwire n_2272 ();
drwire n_2273 ();
drwire n_2274 ();
drwire n_2275 ();
drwire n_2276 ();
drwire n_2277 ();
drwire n_2278 ();
drwire n_2279 ();
drwire n_228 ();
drwire n_2280 ();
drwire n_2281 ();
drwire n_2282 ();
drwire n_2283 ();
drwire n_2284 ();
drwire n_2285 ();
drwire n_2286 ();
drwire n_2287 ();
drwire n_2288 ();
drwire n_2289 ();
drwire n_229 ();
drwire n_2290 ();
drwire n_2291 ();
drwire n_2292 ();
drwire n_2293 ();
drwire n_2294 ();
drwire n_2295 ();
drwire n_2296 ();
drwire n_2297 ();
drwire n_2298 ();
drwire n_2299 ();
drwire n_23 ();
drwire n_230 ();
drwire n_2300 ();
drwire n_2303 ();
drwire n_2304 ();
drwire n_2305 ();
drwire n_2308 ();
drwire n_2309 ();
drwire n_231 ();
drwire n_2310 ();
drwire n_2311 ();
drwire n_2312 ();
drwire n_2313 ();
drwire n_2314 ();
drwire n_2315 ();
drwire n_2316 ();
drwire n_2317 ();
drwire n_2318 ();
drwire n_2319 ();
drwire n_232 ();
drwire n_2320 ();
drwire n_2321 ();
drwire n_2322 ();
drwire n_2323 ();
drwire n_2325 ();
drwire n_2326 ();
drwire n_2327 ();
drwire n_2328 ();
drwire n_2329 ();
drwire n_233 ();
drwire n_2330 ();
drwire n_2331 ();
drwire n_2332 ();
drwire n_2333 ();
drwire n_2334 ();
drwire n_2335 ();
drwire n_2336 ();
drwire n_2337 ();
drwire n_2338 ();
drwire n_2339 ();
drwire n_234 ();
drwire n_2340 ();
drwire n_2341 ();
drwire n_2346 ();
drwire n_2347 ();
drwire n_235 ();
drwire n_2352 ();
drwire n_2353 ();
drwire n_2356 ();
drwire n_236 ();
drwire n_2362 ();
drwire n_2363 ();
drwire n_2364 ();
drwire n_2365 ();
drwire n_2366 ();
drwire n_237 ();
drwire n_2370 ();
drwire n_2373 ();
drwire n_2377 ();
drwire n_2378 ();
drwire n_2379 ();
drwire n_238 ();
drwire n_2380 ();
drwire n_2384 ();
drwire n_2387 ();
drwire n_2388 ();
drwire n_2389 ();
drwire n_239 ();
drwire n_2390 ();
drwire n_2391 ();
drwire n_2392 ();
drwire n_2393 ();
drwire n_2394 ();
drwire n_2395 ();
drwire n_2396 ();
drwire n_2397 ();
drwire n_2399 ();
drwire n_24 ();
drwire n_240 ();
drwire n_2400 ();
drwire n_2401 ();
drwire n_2402 ();
drwire n_2403 ();
drwire n_2404 ();
drwire n_2405 ();
drwire n_2406 ();
drwire n_2407 ();
drwire n_2408 ();
drwire n_2409 ();
drwire n_241 ();
drwire n_2410 ();
drwire n_2411 ();
drwire n_2412 ();
drwire n_2414 ();
drwire n_2415 ();
drwire n_2416 ();
drwire n_2417 ();
drwire n_2418 ();
drwire n_2419 ();
drwire n_242 ();
drwire n_2420 ();
drwire n_2421 ();
drwire n_2422 ();
drwire n_2423 ();
drwire n_2424 ();
drwire n_2425 ();
drwire n_2426 ();
drwire n_2427 ();
drwire n_2428 ();
drwire n_243 ();
drwire n_2430 ();
drwire n_2431 ();
drwire n_2432 ();
drwire n_2433 ();
drwire n_2434 ();
drwire n_2435 ();
drwire n_2436 ();
drwire n_2437 ();
drwire n_2438 ();
drwire n_2439 ();
drwire n_244 ();
drwire n_2440 ();
drwire n_2441 ();
drwire n_2442 ();
drwire n_2443 ();
drwire n_2444 ();
drwire n_2445 ();
drwire n_2446 ();
drwire n_2447 ();
drwire n_2448 ();
drwire n_2449 ();
drwire n_245 ();
drwire n_2450 ();
drwire n_2451 ();
drwire n_2452 ();
drwire n_2453 ();
drwire n_2454 ();
drwire n_2455 ();
drwire n_2456 ();
drwire n_2457 ();
drwire n_2458 ();
drwire n_2459 ();
drwire n_246 ();
drwire n_2460 ();
drwire n_2461 ();
drwire n_2462 ();
drwire n_2463 ();
drwire n_2467 ();
drwire n_247 ();
drwire n_2470 ();
drwire n_2471 ();
drwire n_2472 ();
drwire n_2473 ();
drwire n_2474 ();
drwire n_2475 ();
drwire n_2476 ();
drwire n_2477 ();
drwire n_2478 ();
drwire n_2479 ();
drwire n_248 ();
drwire n_2480 ();
drwire n_2481 ();
drwire n_2482 ();
drwire n_2483 ();
drwire n_2484 ();
drwire n_2485 ();
drwire n_2487 ();
drwire n_2488 ();
drwire n_2489 ();
drwire n_249 ();
drwire n_2490 ();
drwire n_2491 ();
drwire n_2492 ();
drwire n_2493 ();
drwire n_2494 ();
drwire n_2495 ();
drwire n_2496 ();
drwire n_2497 ();
drwire n_2498 ();
drwire n_2499 ();
drwire n_25 ();
drwire n_250 ();
drwire n_2500 ();
drwire n_2502 ();
drwire n_2503 ();
drwire n_2504 ();
drwire n_2505 ();
drwire n_2506 ();
drwire n_2507 ();
drwire n_2509 ();
drwire n_251 ();
drwire n_2510 ();
drwire n_2511 ();
drwire n_2512 ();
drwire n_2513 ();
drwire n_2515 ();
drwire n_2516 ();
drwire n_2517 ();
drwire n_2518 ();
drwire n_2519 ();
drwire n_252 ();
drwire n_2520 ();
drwire n_2523 ();
drwire n_2526 ();
drwire n_253 ();
drwire n_2531 ();
drwire n_2534 ();
drwire n_2535 ();
drwire n_2536 ();
drwire n_254 ();
drwire n_2541 ();
drwire n_2542 ();
drwire n_2543 ();
drwire n_2544 ();
drwire n_2545 ();
drwire n_2546 ();
drwire n_2547 ();
drwire n_2548 ();
drwire n_2549 ();
drwire n_255 ();
drwire n_2550 ();
drwire n_2551 ();
drwire n_2552 ();
drwire n_2553 ();
drwire n_2554 ();
drwire n_2555 ();
drwire n_2556 ();
drwire n_2557 ();
drwire n_2558 ();
drwire n_2559 ();
drwire n_256 ();
drwire n_2560 ();
drwire n_2561 ();
drwire n_2562 ();
drwire n_2563 ();
drwire n_2564 ();
drwire n_2565 ();
drwire n_2566 ();
drwire n_2568 ();
drwire n_2569 ();
drwire n_257 ();
drwire n_2570 ();
drwire n_2571 ();
drwire n_2572 ();
drwire n_2573 ();
drwire n_2574 ();
drwire n_2575 ();
drwire n_2576 ();
drwire n_2577 ();
drwire n_2578 ();
drwire n_2579 ();
drwire n_258 ();
drwire n_2580 ();
drwire n_2581 ();
drwire n_2582 ();
drwire n_2583 ();
drwire n_2584 ();
drwire n_2585 ();
drwire n_2586 ();
drwire n_2587 ();
drwire n_2588 ();
drwire n_2589 ();
drwire n_259 ();
drwire n_2590 ();
drwire n_2591 ();
drwire n_2592 ();
drwire n_2593 ();
drwire n_2594 ();
drwire n_2595 ();
drwire n_2596 ();
drwire n_2597 ();
drwire n_2598 ();
drwire n_2599 ();
drwire n_26 ();
drwire n_260 ();
drwire n_2600 ();
drwire n_2601 ();
drwire n_2602 ();
drwire n_261 ();
drwire n_2610 ();
drwire n_2612 ();
drwire n_2614 ();
drwire n_2615 ();
drwire n_2616 ();
drwire n_2617 ();
drwire n_2618 ();
drwire n_2619 ();
drwire n_262 ();
drwire n_2624 ();
drwire n_2625 ();
drwire n_2626 ();
drwire n_2627 ();
drwire n_2628 ();
drwire n_2629 ();
drwire n_263 ();
drwire n_2630 ();
drwire n_2633 ();
drwire n_2634 ();
drwire n_2636 ();
drwire n_2637 ();
drwire n_2638 ();
drwire n_264 ();
drwire n_2640 ();
drwire n_2641 ();
drwire n_2642 ();
drwire n_2644 ();
drwire n_2645 ();
drwire n_2646 ();
drwire n_2647 ();
drwire n_2648 ();
drwire n_2649 ();
drwire n_265 ();
drwire n_2650 ();
drwire n_2651 ();
drwire n_2652 ();
drwire n_2653 ();
drwire n_2654 ();
drwire n_2656 ();
drwire n_2657 ();
drwire n_2658 ();
drwire n_2659 ();
drwire n_266 ();
drwire n_2660 ();
drwire n_2661 ();
drwire n_2662 ();
drwire n_2663 ();
drwire n_2664 ();
drwire n_2665 ();
drwire n_2666 ();
drwire n_2667 ();
drwire n_2669 ();
drwire n_267 ();
drwire n_2670 ();
drwire n_2671 ();
drwire n_2673 ();
drwire n_2674 ();
drwire n_2675 ();
drwire n_2679 ();
drwire n_268 ();
drwire n_2680 ();
drwire n_2681 ();
drwire n_2682 ();
drwire n_2683 ();
drwire n_2686 ();
drwire n_2687 ();
drwire n_2688 ();
drwire n_2689 ();
drwire n_269 ();
drwire n_2690 ();
drwire n_2692 ();
drwire n_2693 ();
drwire n_2696 ();
drwire n_27 ();
drwire n_270 ();
drwire n_2702 ();
drwire n_2704 ();
drwire n_2705 ();
drwire n_2708 ();
drwire n_2709 ();
drwire n_271 ();
drwire n_2711 ();
drwire n_2712 ();
drwire n_2713 ();
drwire n_2714 ();
drwire n_2715 ();
drwire n_2716 ();
drwire n_2717 ();
drwire n_2718 ();
drwire n_2719 ();
drwire n_272 ();
drwire n_2720 ();
drwire n_2724 ();
drwire n_2725 ();
drwire n_2726 ();
drwire n_2728 ();
drwire n_2729 ();
drwire n_273 ();
drwire n_2730 ();
drwire n_2731 ();
drwire n_2732 ();
drwire n_2733 ();
drwire n_2734 ();
drwire n_2735 ();
drwire n_2736 ();
drwire n_2737 ();
drwire n_2738 ();
drwire n_2739 ();
drwire n_274 ();
drwire n_2740 ();
drwire n_2741 ();
drwire n_2743 ();
drwire n_2749 ();
drwire n_275 ();
drwire n_2750 ();
drwire n_2753 ();
drwire n_2755 ();
drwire n_2756 ();
drwire n_2757 ();
drwire n_2758 ();
drwire n_2759 ();
drwire n_276 ();
drwire n_2760 ();
drwire n_2761 ();
drwire n_2762 ();
drwire n_2763 ();
drwire n_2764 ();
drwire n_2765 ();
drwire n_2766 ();
drwire n_2769 ();
drwire n_277 ();
drwire n_2770 ();
drwire n_2771 ();
drwire n_2772 ();
drwire n_278 ();
drwire n_279 ();
drwire n_2792 ();
drwire n_2793 ();
drwire n_2798 ();
drwire n_28 ();
drwire n_280 ();
drwire n_2805 ();
drwire n_2807 ();
drwire n_281 ();
drwire n_2812 ();
drwire n_2813 ();
drwire n_2814 ();
drwire n_2815 ();
drwire n_2816 ();
drwire n_2817 ();
drwire n_2818 ();
drwire n_2819 ();
drwire n_282 ();
drwire n_2820 ();
drwire n_2821 ();
drwire n_2823 ();
drwire n_2824 ();
drwire n_2825 ();
drwire n_2826 ();
drwire n_2827 ();
drwire n_2828 ();
drwire n_283 ();
drwire n_2831 ();
drwire n_2832 ();
drwire n_2833 ();
drwire n_284 ();
drwire n_2841 ();
drwire n_2842 ();
drwire n_2843 ();
drwire n_2846 ();
drwire n_285 ();
drwire n_2852 ();
drwire n_2853 ();
drwire n_2854 ();
drwire n_286 ();
drwire n_2862 ();
drwire n_2866 ();
drwire n_2867 ();
drwire n_2868 ();
drwire n_2869 ();
drwire n_287 ();
drwire n_2870 ();
drwire n_2871 ();
drwire n_2872 ();
drwire n_2873 ();
drwire n_2874 ();
drwire n_2875 ();
drwire n_2876 ();
drwire n_2877 ();
drwire n_2878 ();
drwire n_2879 ();
drwire n_288 ();
drwire n_2880 ();
drwire n_2881 ();
drwire n_289 ();
drwire n_29 ();
drwire n_290 ();
drwire n_2901 ();
drwire n_2902 ();
drwire n_2903 ();
drwire n_2904 ();
drwire n_2905 ();
drwire n_2909 ();
drwire n_291 ();
drwire n_2910 ();
drwire n_2911 ();
drwire n_2912 ();
drwire n_2914 ();
drwire n_2915 ();
drwire n_2916 ();
drwire n_2917 ();
drwire n_2918 ();
drwire n_2919 ();
drwire n_292 ();
drwire n_2920 ();
drwire n_2921 ();
drwire n_2922 ();
drwire n_2923 ();
drwire n_2924 ();
drwire n_2925 ();
drwire n_2926 ();
drwire n_2927 ();
drwire n_2928 ();
drwire n_2929 ();
drwire n_293 ();
drwire n_2931 ();
drwire n_2932 ();
drwire n_2933 ();
drwire n_2934 ();
drwire n_2935 ();
drwire n_2937 ();
drwire n_2938 ();
drwire n_2939 ();
drwire n_294 ();
drwire n_2940 ();
drwire n_2941 ();
drwire n_2942 ();
drwire n_2943 ();
drwire n_2944 ();
drwire n_2945 ();
drwire n_2946 ();
drwire n_2947 ();
drwire n_2949 ();
drwire n_295 ();
drwire n_2950 ();
drwire n_2952 ();
drwire n_2953 ();
drwire n_2954 ();
drwire n_2955 ();
drwire n_2956 ();
drwire n_2958 ();
drwire n_2959 ();
drwire n_296 ();
drwire n_2960 ();
drwire n_2961 ();
drwire n_2963 ();
drwire n_2966 ();
drwire n_297 ();
drwire n_298 ();
drwire n_2981 ();
drwire n_2982 ();
drwire n_2983 ();
drwire n_299 ();
drwire n_2993 ();
drwire n_2994 ();
drwire n_2995 ();
drwire n_2996 ();
drwire n_2997 ();
drwire n_2998 ();
drwire n_3 ();
drwire n_30 ();
drwire n_300 ();
drwire n_3008 ();
drwire n_301 ();
drwire n_3010 ();
drwire n_3011 ();
drwire n_302 ();
drwire n_303 ();
drwire n_304 ();
drwire n_305 ();
drwire n_306 ();
drwire n_307 ();
drwire n_308 ();
drwire n_309 ();
drwire n_31 ();
drwire n_310 ();
drwire n_3109 ();
drwire n_311 ();
drwire n_3110 ();
drwire n_3111 ();
drwire n_3112 ();
drwire n_312 ();
drwire n_3125 ();
drwire n_3126 ();
drwire n_3127 ();
drwire n_3128 ();
drwire n_3129 ();
drwire n_313 ();
drwire n_3130 ();
drwire n_3131 ();
drwire n_3134 ();
drwire n_3139 ();
drwire n_314 ();
drwire n_3141 ();
drwire n_3142 ();
drwire n_3143 ();
drwire n_3144 ();
drwire n_3145 ();
drwire n_315 ();
drwire n_3157 ();
drwire n_3158 ();
drwire n_3159 ();
drwire n_316 ();
drwire n_3160 ();
drwire n_3161 ();
drwire n_3162 ();
drwire n_3163 ();
drwire n_3164 ();
drwire n_3165 ();
drwire n_3166 ();
drwire n_3167 ();
drwire n_3168 ();
drwire n_3169 ();
drwire n_317 ();
drwire n_3170 ();
drwire n_3172 ();
drwire n_3177 ();
drwire n_3179 ();
drwire n_318 ();
drwire n_3180 ();
drwire n_3181 ();
drwire n_3182 ();
drwire n_3183 ();
drwire n_3184 ();
drwire n_3185 ();
drwire n_3186 ();
drwire n_3187 ();
drwire n_3188 ();
drwire n_3189 ();
drwire n_319 ();
drwire n_3190 ();
drwire n_3191 ();
drwire n_3192 ();
drwire n_3194 ();
drwire n_3199 ();
drwire n_32 ();
drwire n_320 ();
drwire n_3201 ();
drwire n_3202 ();
drwire n_3203 ();
drwire n_3204 ();
drwire n_3207 ();
drwire n_3209 ();
drwire n_321 ();
drwire n_3214 ();
drwire n_3217 ();
drwire n_322 ();
drwire n_3222 ();
drwire n_3225 ();
drwire n_323 ();
drwire n_3230 ();
drwire n_3232 ();
drwire n_3233 ();
drwire n_3236 ();
drwire n_3237 ();
drwire n_3239 ();
drwire n_324 ();
drwire n_3244 ();
drwire n_3247 ();
drwire n_325 ();
drwire n_3252 ();
drwire n_3255 ();
drwire n_326 ();
drwire n_3260 ();
drwire n_3262 ();
drwire n_3263 ();
drwire n_3264 ();
drwire n_3265 ();
drwire n_3268 ();
drwire n_3269 ();
drwire n_327 ();
drwire n_3270 ();
drwire n_3271 ();
drwire n_3272 ();
drwire n_3273 ();
drwire n_3274 ();
drwire n_3275 ();
drwire n_3276 ();
drwire n_3277 ();
drwire n_3278 ();
drwire n_3279 ();
drwire n_328 ();
drwire n_3283 ();
drwire n_3284 ();
drwire n_3289 ();
drwire n_329 ();
drwire n_3290 ();
drwire n_3291 ();
drwire n_3292 ();
drwire n_3293 ();
drwire n_3294 ();
drwire n_3296 ();
drwire n_3297 ();
drwire n_3298 ();
drwire n_3299 ();
drwire n_33 ();
drwire n_330 ();
drwire n_3300 ();
drwire n_331 ();
drwire n_3311 ();
drwire n_3315 ();
drwire n_3316 ();
drwire n_3317 ();
drwire n_3318 ();
drwire n_3319 ();
drwire n_332 ();
drwire n_3320 ();
drwire n_3321 ();
drwire n_3322 ();
drwire n_3323 ();
drwire n_3324 ();
drwire n_3325 ();
drwire n_3326 ();
drwire n_3327 ();
drwire n_3328 ();
drwire n_3329 ();
drwire n_333 ();
drwire n_3330 ();
drwire n_3331 ();
drwire n_3332 ();
drwire n_3333 ();
drwire n_3334 ();
drwire n_3335 ();
drwire n_3336 ();
drwire n_3337 ();
drwire n_3338 ();
drwire n_3339 ();
drwire n_334 ();
drwire n_3340 ();
drwire n_3341 ();
drwire n_3342 ();
drwire n_3343 ();
drwire n_3344 ();
drwire n_3345 ();
drwire n_3346 ();
drwire n_3347 ();
drwire n_3348 ();
drwire n_3349 ();
drwire n_335 ();
drwire n_3350 ();
drwire n_3351 ();
drwire n_3352 ();
drwire n_3353 ();
drwire n_3355 ();
drwire n_3356 ();
drwire n_3357 ();
drwire n_3358 ();
drwire n_3359 ();
drwire n_336 ();
drwire n_3360 ();
drwire n_3361 ();
drwire n_3362 ();
drwire n_3363 ();
drwire n_3364 ();
drwire n_3365 ();
drwire n_3366 ();
drwire n_3367 ();
drwire n_3368 ();
drwire n_3369 ();
drwire n_337 ();
drwire n_3370 ();
drwire n_3371 ();
drwire n_3372 ();
drwire n_3375 ();
drwire n_3376 ();
drwire n_3377 ();
drwire n_3378 ();
drwire n_3379 ();
drwire n_338 ();
drwire n_3380 ();
drwire n_339 ();
drwire n_3399 ();
drwire n_340 ();
drwire n_3400 ();
drwire n_3401 ();
drwire n_3402 ();
drwire n_3403 ();
drwire n_3404 ();
drwire n_3405 ();
drwire n_341 ();
drwire n_3418 ();
drwire n_3419 ();
drwire n_342 ();
drwire n_3420 ();
drwire n_3421 ();
drwire n_3422 ();
drwire n_3423 ();
drwire n_3424 ();
drwire n_343 ();
drwire n_3434 ();
drwire n_3435 ();
drwire n_3436 ();
drwire n_3437 ();
drwire n_3438 ();
drwire n_3439 ();
drwire n_344 ();
drwire n_3440 ();
drwire n_3441 ();
drwire n_3442 ();
drwire n_3443 ();
drwire n_3444 ();
drwire n_345 ();
drwire n_3451 ();
drwire n_3452 ();
drwire n_3453 ();
drwire n_3454 ();
drwire n_346 ();
drwire n_347 ();
drwire n_348 ();
drwire n_3487 ();
drwire n_3488 ();
drwire n_3489 ();
drwire n_349 ();
drwire n_3490 ();
drwire n_3491 ();
drwire n_3493 ();
drwire n_35 ();
drwire n_350 ();
drwire n_3502 ();
drwire n_3503 ();
drwire n_3504 ();
drwire n_3505 ();
drwire n_351 ();
drwire n_3514 ();
drwire n_3518 ();
drwire n_3519 ();
drwire n_352 ();
drwire n_3520 ();
drwire n_3521 ();
drwire n_3522 ();
drwire n_3523 ();
drwire n_3524 ();
drwire n_3525 ();
drwire n_3527 ();
drwire n_353 ();
drwire n_355 ();
drwire n_357 ();
drwire n_3571 ();
drwire n_3572 ();
drwire n_3573 ();
drwire n_3574 ();
drwire n_3575 ();
drwire n_3576 ();
drwire n_3577 ();
drwire n_3578 ();
drwire n_3579 ();
drwire n_358 ();
drwire n_3580 ();
drwire n_359 ();
drwire n_3591 ();
drwire n_3592 ();
drwire n_3593 ();
drwire n_3594 ();
drwire n_3595 ();
drwire n_3596 ();
drwire n_3597 ();
drwire n_3598 ();
drwire n_3599 ();
drwire n_36 ();
drwire n_360 ();
drwire n_3600 ();
drwire n_3607 ();
drwire n_3609 ();
drwire n_361 ();
drwire n_3611 ();
drwire n_3612 ();
drwire n_3613 ();
drwire n_3614 ();
drwire n_3615 ();
drwire n_3616 ();
drwire n_3618 ();
drwire n_3619 ();
drwire n_362 ();
drwire n_3624 ();
drwire n_3625 ();
drwire n_3626 ();
drwire n_3627 ();
drwire n_3628 ();
drwire n_3629 ();
drwire n_363 ();
drwire n_3630 ();
drwire n_3631 ();
drwire n_3632 ();
drwire n_3633 ();
drwire n_3634 ();
drwire n_3635 ();
drwire n_3636 ();
drwire n_3637 ();
drwire n_3638 ();
drwire n_364 ();
drwire n_3640 ();
drwire n_3641 ();
drwire n_3643 ();
drwire n_3644 ();
drwire n_3645 ();
drwire n_3646 ();
drwire n_3648 ();
drwire n_3649 ();
drwire n_365 ();
drwire n_3650 ();
drwire n_3651 ();
drwire n_3652 ();
drwire n_3655 ();
drwire n_3656 ();
drwire n_3657 ();
drwire n_3658 ();
drwire n_3659 ();
drwire n_366 ();
drwire n_3660 ();
drwire n_3661 ();
drwire n_3662 ();
drwire n_3663 ();
drwire n_3664 ();
drwire n_3667 ();
drwire n_3668 ();
drwire n_367 ();
drwire n_3671 ();
drwire n_3677 ();
drwire n_3678 ();
drwire n_3679 ();
drwire n_368 ();
drwire n_3680 ();
drwire n_3681 ();
drwire n_3687 ();
drwire n_3688 ();
drwire n_3689 ();
drwire n_369 ();
drwire n_3690 ();
drwire n_3691 ();
drwire n_3692 ();
drwire n_3693 ();
drwire n_3694 ();
drwire n_3699 ();
drwire n_37 ();
drwire n_370 ();
drwire n_3700 ();
drwire n_3701 ();
drwire n_3702 ();
drwire n_3703 ();
drwire n_3704 ();
drwire n_3705 ();
drwire n_3706 ();
drwire n_3707 ();
drwire n_3708 ();
drwire n_3709 ();
drwire n_371 ();
drwire n_3710 ();
drwire n_3711 ();
drwire n_3712 ();
drwire n_3713 ();
drwire n_3714 ();
drwire n_3715 ();
drwire n_3716 ();
drwire n_3717 ();
drwire n_3718 ();
drwire n_3719 ();
drwire n_372 ();
drwire n_3720 ();
drwire n_3721 ();
drwire n_3722 ();
drwire n_3723 ();
drwire n_3724 ();
drwire n_3725 ();
drwire n_3726 ();
drwire n_3727 ();
drwire n_3728 ();
drwire n_3729 ();
drwire n_373 ();
drwire n_3731 ();
drwire n_3732 ();
drwire n_3733 ();
drwire n_3734 ();
drwire n_3735 ();
drwire n_3737 ();
drwire n_3738 ();
drwire n_374 ();
drwire n_3742 ();
drwire n_3743 ();
drwire n_3744 ();
drwire n_375 ();
drwire n_3751 ();
drwire n_3757 ();
drwire n_3758 ();
drwire n_3759 ();
drwire n_376 ();
drwire n_3760 ();
drwire n_3761 ();
drwire n_3764 ();
drwire n_3768 ();
drwire n_377 ();
drwire n_3770 ();
drwire n_3771 ();
drwire n_3777 ();
drwire n_3778 ();
drwire n_3779 ();
drwire n_378 ();
drwire n_379 ();
drwire n_3790 ();
drwire n_3791 ();
drwire n_3792 ();
drwire n_3794 ();
drwire n_3795 ();
drwire n_3796 ();
drwire n_38 ();
drwire n_380 ();
drwire n_3804 ();
drwire n_3805 ();
drwire n_381 ();
drwire n_3813 ();
drwire n_3814 ();
drwire n_3816 ();
drwire n_3817 ();
drwire n_3818 ();
drwire n_3819 ();
drwire n_382 ();
drwire n_3821 ();
drwire n_3825 ();
drwire n_3826 ();
drwire n_3827 ();
drwire n_3828 ();
drwire n_383 ();
drwire n_3830 ();
drwire n_3831 ();
drwire n_3832 ();
drwire n_3833 ();
drwire n_3834 ();
drwire n_3835 ();
drwire n_3836 ();
drwire n_3837 ();
drwire n_3838 ();
drwire n_3839 ();
drwire n_384 ();
drwire n_3840 ();
drwire n_3841 ();
drwire n_3842 ();
drwire n_3843 ();
drwire n_3844 ();
drwire n_3845 ();
drwire n_3847 ();
drwire n_3848 ();
drwire n_3849 ();
drwire n_385 ();
drwire n_3850 ();
drwire n_3851 ();
drwire n_3852 ();
drwire n_3853 ();
drwire n_3854 ();
drwire n_386 ();
drwire n_3861 ();
drwire n_3866 ();
drwire n_3869 ();
drwire n_387 ();
drwire n_3871 ();
drwire n_3872 ();
drwire n_3874 ();
drwire n_3875 ();
drwire n_3876 ();
drwire n_3877 ();
drwire n_3878 ();
drwire n_3879 ();
drwire n_388 ();
drwire n_3880 ();
drwire n_3881 ();
drwire n_3886 ();
drwire n_3887 ();
drwire n_3888 ();
drwire n_389 ();
drwire n_3890 ();
drwire n_3891 ();
drwire n_3892 ();
drwire n_3893 ();
drwire n_3894 ();
drwire n_3895 ();
drwire n_3896 ();
drwire n_39 ();
drwire n_390 ();
drwire n_3900 ();
drwire n_3901 ();
drwire n_3902 ();
drwire n_3903 ();
drwire n_3904 ();
drwire n_3905 ();
drwire n_3906 ();
drwire n_3907 ();
drwire n_3908 ();
drwire n_3909 ();
drwire n_391 ();
drwire n_3910 ();
drwire n_3911 ();
drwire n_3912 ();
drwire n_3913 ();
drwire n_3914 ();
drwire n_392 ();
drwire n_3926 ();
drwire n_3927 ();
drwire n_3928 ();
drwire n_393 ();
drwire n_3930 ();
drwire n_3931 ();
drwire n_3932 ();
drwire n_3933 ();
drwire n_3934 ();
drwire n_3935 ();
drwire n_3936 ();
drwire n_394 ();
drwire n_3941 ();
drwire n_3942 ();
drwire n_3943 ();
drwire n_3944 ();
drwire n_3945 ();
drwire n_3946 ();
drwire n_3947 ();
drwire n_3948 ();
drwire n_3949 ();
drwire n_395 ();
drwire n_3950 ();
drwire n_3951 ();
drwire n_3952 ();
drwire n_3953 ();
drwire n_3954 ();
drwire n_3955 ();
drwire n_3956 ();
drwire n_3958 ();
drwire n_3959 ();
drwire n_396 ();
drwire n_3960 ();
drwire n_3961 ();
drwire n_3962 ();
drwire n_3963 ();
drwire n_3964 ();
drwire n_3965 ();
drwire n_3966 ();
drwire n_3967 ();
drwire n_3968 ();
drwire n_3969 ();
drwire n_397 ();
drwire n_3970 ();
drwire n_3972 ();
drwire n_3973 ();
drwire n_3974 ();
drwire n_3975 ();
drwire n_3976 ();
drwire n_3977 ();
drwire n_3978 ();
drwire n_3979 ();
drwire n_398 ();
drwire n_3980 ();
drwire n_3981 ();
drwire n_3982 ();
drwire n_3983 ();
drwire n_3984 ();
drwire n_3985 ();
drwire n_3986 ();
drwire n_3988 ();
drwire n_3989 ();
drwire n_399 ();
drwire n_3997 ();
drwire n_3998 ();
drwire n_3999 ();
drwire n_4 ();
drwire n_40 ();
drwire n_400 ();
drwire n_4000 ();
drwire n_4001 ();
drwire n_4002 ();
drwire n_4003 ();
drwire n_401 ();
drwire n_4017 ();
drwire n_4018 ();
drwire n_4019 ();
drwire n_402 ();
drwire n_4020 ();
drwire n_4021 ();
drwire n_4022 ();
drwire n_4023 ();
drwire n_4024 ();
drwire n_4025 ();
drwire n_4026 ();
drwire n_4027 ();
drwire n_4028 ();
drwire n_4029 ();
drwire n_403 ();
drwire n_4030 ();
drwire n_4031 ();
drwire n_404 ();
drwire n_4046 ();
drwire n_4048 ();
drwire n_4049 ();
drwire n_405 ();
drwire n_4055 ();
drwire n_4057 ();
drwire n_4058 ();
drwire n_4059 ();
drwire n_406 ();
drwire n_4060 ();
drwire n_4061 ();
drwire n_4062 ();
drwire n_407 ();
drwire n_408 ();
drwire n_4087 ();
drwire n_4088 ();
drwire n_4089 ();
drwire n_409 ();
drwire n_4090 ();
drwire n_4091 ();
drwire n_4092 ();
drwire n_4099 ();
drwire n_410 ();
drwire n_4100 ();
drwire n_411 ();
drwire n_412 ();
drwire n_413 ();
drwire n_4135 ();
drwire n_4136 ();
drwire n_4137 ();
drwire n_4138 ();
drwire n_414 ();
drwire n_415 ();
drwire n_416 ();
drwire n_417 ();
drwire n_418 ();
drwire n_419 ();
drwire n_42 ();
drwire n_420 ();
drwire n_421 ();
drwire n_422 ();
drwire n_423 ();
drwire n_424 ();
drwire n_425 ();
drwire n_4257 ();
drwire n_4258 ();
drwire n_4259 ();
drwire n_426 ();
drwire n_427 ();
drwire n_4277 ();
drwire n_4278 ();
drwire n_4279 ();
drwire n_428 ();
drwire n_4280 ();
drwire n_4281 ();
drwire n_4282 ();
drwire n_4283 ();
drwire n_4289 ();
drwire n_429 ();
drwire n_4290 ();
drwire n_4291 ();
drwire n_4292 ();
drwire n_4293 ();
drwire n_4294 ();
drwire n_4295 ();
drwire n_4296 ();
drwire n_4297 ();
drwire n_4298 ();
drwire n_4299 ();
drwire n_43 ();
drwire n_430 ();
drwire n_4300 ();
drwire n_4301 ();
drwire n_4302 ();
drwire n_4303 ();
drwire n_4304 ();
drwire n_4305 ();
drwire n_4306 ();
drwire n_431 ();
drwire n_432 ();
drwire n_433 ();
drwire n_4331 ();
drwire n_4332 ();
drwire n_4334 ();
drwire n_4335 ();
drwire n_4336 ();
drwire n_4337 ();
drwire n_434 ();
drwire n_435 ();
drwire n_4350 ();
drwire n_4351 ();
drwire n_4352 ();
drwire n_4353 ();
drwire n_4354 ();
drwire n_4355 ();
drwire n_4356 ();
drwire n_4358 ();
drwire n_436 ();
drwire n_4363 ();
drwire n_4365 ();
drwire n_4366 ();
drwire n_4367 ();
drwire n_4368 ();
drwire n_4369 ();
drwire n_437 ();
drwire n_4370 ();
drwire n_4371 ();
drwire n_4372 ();
drwire n_4377 ();
drwire n_438 ();
drwire n_4380 ();
drwire n_439 ();
drwire n_4397 ();
drwire n_4398 ();
drwire n_4399 ();
drwire n_44 ();
drwire n_440 ();
drwire n_4400 ();
drwire n_4401 ();
drwire n_4402 ();
drwire n_4403 ();
drwire n_4404 ();
drwire n_4405 ();
drwire n_4406 ();
drwire n_4407 ();
drwire n_4408 ();
drwire n_4409 ();
drwire n_441 ();
drwire n_4410 ();
drwire n_4411 ();
drwire n_442 ();
drwire n_443 ();
drwire n_444 ();
drwire n_445 ();
drwire n_446 ();
drwire n_447 ();
drwire n_448 ();
drwire n_449 ();
drwire n_4498 ();
drwire n_4499 ();
drwire n_45 ();
drwire n_450 ();
drwire n_4500 ();
drwire n_4501 ();
drwire n_4502 ();
drwire n_452 ();
drwire n_4549 ();
drwire n_455 ();
drwire n_4550 ();
drwire n_4552 ();
drwire n_4557 ();
drwire n_4558 ();
drwire n_457 ();
drwire n_459 ();
drwire n_4597 ();
drwire n_46 ();
drwire n_460 ();
drwire n_461 ();
drwire n_462 ();
drwire n_463 ();
drwire n_464 ();
drwire n_465 ();
drwire n_466 ();
drwire n_467 ();
drwire n_468 ();
drwire n_469 ();
drwire n_47 ();
drwire n_470 ();
drwire n_471 ();
drwire n_472 ();
drwire n_473 ();
drwire n_474 ();
drwire n_475 ();
drwire n_476 ();
drwire n_477 ();
drwire n_478 ();
drwire n_479 ();
drwire n_48 ();
drwire n_480 ();
drwire n_481 ();
drwire n_482 ();
drwire n_483 ();
drwire n_484 ();
drwire n_485 ();
drwire n_486 ();
drwire n_487 ();
drwire n_488 ();
drwire n_489 ();
drwire n_49 ();
drwire n_490 ();
drwire n_491 ();
drwire n_492 ();
drwire n_493 ();
drwire n_494 ();
drwire n_495 ();
drwire n_496 ();
drwire n_497 ();
drwire n_5 ();
drwire n_50 ();
drwire n_500 ();
drwire n_501 ();
drwire n_502 ();
drwire n_503 ();
drwire n_504 ();
drwire n_505 ();
drwire n_506 ();
drwire n_507 ();
drwire n_508 ();
drwire n_509 ();
drwire n_51 ();
drwire n_510 ();
drwire n_511 ();
drwire n_512 ();
drwire n_514 ();
drwire n_515 ();
drwire n_516 ();
drwire n_517 ();
drwire n_518 ();
drwire n_519 ();
drwire n_52 ();
drwire n_520 ();
drwire n_521 ();
drwire n_522 ();
drwire n_523 ();
drwire n_524 ();
drwire n_525 ();
drwire n_526 ();
drwire n_527 ();
drwire n_528 ();
drwire n_529 ();
drwire n_53 ();
drwire n_530 ();
drwire n_531 ();
drwire n_532 ();
drwire n_533 ();
drwire n_534 ();
drwire n_535 ();
drwire n_536 ();
drwire n_537 ();
drwire n_538 ();
drwire n_539 ();
drwire n_54 ();
drwire n_540 ();
drwire n_541 ();
drwire n_542 ();
drwire n_543 ();
drwire n_544 ();
drwire n_545 ();
drwire n_546 ();
drwire n_547 ();
drwire n_548 ();
drwire n_549 ();
drwire n_55 ();
drwire n_550 ();
drwire n_551 ();
drwire n_552 ();
drwire n_553 ();
drwire n_554 ();
drwire n_555 ();
drwire n_556 ();
drwire n_557 ();
drwire n_558 ();
drwire n_559 ();
drwire n_56 ();
drwire n_560 ();
drwire n_561 ();
drwire n_562 ();
drwire n_563 ();
drwire n_564 ();
drwire n_565 ();
drwire n_566 ();
drwire n_567 ();
drwire n_568 ();
drwire n_569 ();
drwire n_57 ();
drwire n_570 ();
drwire n_571 ();
drwire n_572 ();
drwire n_573 ();
drwire n_574 ();
drwire n_575 ();
drwire n_576 ();
drwire n_577 ();
drwire n_578 ();
drwire n_579 ();
drwire n_58 ();
drwire n_581 ();
drwire n_584 ();
drwire n_585 ();
drwire n_586 ();
drwire n_587 ();
drwire n_588 ();
drwire n_589 ();
drwire n_59 ();
drwire n_590 ();
drwire n_591 ();
drwire n_592 ();
drwire n_593 ();
drwire n_594 ();
drwire n_595 ();
drwire n_596 ();
drwire n_597 ();
drwire n_598 ();
drwire n_599 ();
drwire n_6 ();
drwire n_60 ();
drwire n_603 ();
drwire n_604 ();
drwire n_606 ();
drwire n_607 ();
drwire n_608 ();
drwire n_609 ();
drwire n_61 ();
drwire n_610 ();
drwire n_611 ();
drwire n_612 ();
drwire n_613 ();
drwire n_614 ();
drwire n_615 ();
drwire n_616 ();
drwire n_617 ();
drwire n_618 ();
drwire n_619 ();
drwire n_62 ();
drwire n_620 ();
drwire n_621 ();
drwire n_622 ();
drwire n_623 ();
drwire n_624 ();
drwire n_625 ();
drwire n_626 ();
drwire n_627 ();
drwire n_628 ();
drwire n_629 ();
drwire n_63 ();
drwire n_630 ();
drwire n_631 ();
drwire n_632 ();
drwire n_633 ();
drwire n_634 ();
drwire n_635 ();
drwire n_636 ();
drwire n_637 ();
drwire n_638 ();
drwire n_639 ();
drwire n_64 ();
drwire n_640 ();
drwire n_641 ();
drwire n_642 ();
drwire n_643 ();
drwire n_644 ();
drwire n_645 ();
drwire n_646 ();
drwire n_647 ();
drwire n_648 ();
drwire n_649 ();
drwire n_65 ();
drwire n_650 ();
drwire n_652 ();
drwire n_653 ();
drwire n_654 ();
drwire n_655 ();
drwire n_659 ();
drwire n_66 ();
drwire n_660 ();
drwire n_661 ();
drwire n_662 ();
drwire n_663 ();
drwire n_664 ();
drwire n_665 ();
drwire n_666 ();
drwire n_667 ();
drwire n_668 ();
drwire n_669 ();
drwire n_67 ();
drwire n_670 ();
drwire n_671 ();
drwire n_672 ();
drwire n_673 ();
drwire n_674 ();
drwire n_675 ();
drwire n_676 ();
drwire n_677 ();
drwire n_678 ();
drwire n_679 ();
drwire n_68 ();
drwire n_680 ();
drwire n_681 ();
drwire n_682 ();
drwire n_683 ();
drwire n_684 ();
drwire n_685 ();
drwire n_686 ();
drwire n_687 ();
drwire n_688 ();
drwire n_69 ();
drwire n_693 ();
drwire n_694 ();
drwire n_695 ();
drwire n_696 ();
drwire n_697 ();
drwire n_698 ();
drwire n_699 ();
drwire n_7 ();
drwire n_70 ();
drwire n_700 ();
drwire n_701 ();
drwire n_702 ();
drwire n_703 ();
drwire n_704 ();
drwire n_705 ();
drwire n_706 ();
drwire n_707 ();
drwire n_708 ();
drwire n_709 ();
drwire n_71 ();
drwire n_710 ();
drwire n_711 ();
drwire n_712 ();
drwire n_713 ();
drwire n_714 ();
drwire n_715 ();
drwire n_716 ();
drwire n_717 ();
drwire n_718 ();
drwire n_719 ();
drwire n_72 ();
drwire n_721 ();
drwire n_722 ();
drwire n_724 ();
drwire n_728 ();
drwire n_73 ();
drwire n_736 ();
drwire n_74 ();
drwire n_75 ();
drwire n_76 ();
drwire n_764 ();
drwire n_765 ();
drwire n_766 ();
drwire n_77 ();
drwire n_776 ();
drwire n_777 ();
drwire n_778 ();
drwire n_78 ();
drwire n_788 ();
drwire n_789 ();
drwire n_79 ();
drwire n_790 ();
drwire n_794 ();
drwire n_795 ();
drwire n_796 ();
drwire n_797 ();
drwire n_798 ();
drwire n_799 ();
drwire n_8 ();
drwire n_80 ();
drwire n_801 ();
drwire n_81 ();
drwire n_82 ();
drwire n_825 ();
drwire n_83 ();
drwire n_84 ();
drwire n_848 ();
drwire n_849 ();
drwire n_85 ();
drwire n_850 ();
drwire n_86 ();
drwire n_87 ();
drwire n_874 ();
drwire n_88 ();
drwire n_89 ();
drwire n_9 ();
drwire n_90 ();
drwire n_91 ();
drwire n_92 ();
drwire n_93 ();
drwire n_938 ();
drwire n_939 ();
drwire n_94 ();
drwire n_940 ();
drwire n_941 ();
drwire n_942 ();
drwire n_943 ();
drwire n_944 ();
drwire n_945 ();
drwire n_946 ();
drwire n_947 ();
drwire n_948 ();
drwire n_949 ();
drwire n_95 ();
drwire n_950 ();
drwire n_951 ();
drwire n_952 ();
drwire n_953 ();
drwire n_954 ();
drwire n_955 ();
drwire n_956 ();
drwire n_957 ();
drwire n_958 ();
drwire n_959 ();
drwire n_96 ();
drwire n_960 ();
drwire n_961 ();
drwire n_962 ();
drwire n_963 ();
drwire n_964 ();
drwire n_965 ();
drwire n_966 ();
drwire n_967 ();
drwire n_968 ();
drwire n_97 ();
drwire n_974 ();
drwire n_975 ();
drwire n_98 ();
drwire n_981 ();
drwire n_983 ();
drwire n_985 ();
drwire n_986 ();
drwire n_987 ();
drwire n_988 ();
drwire n_99 ();
drwire ps_0_ ();
drwire ps_1_ ();
drwire sum_0_ ();
drwire sum_10_ ();
drwire sum_11_ ();
drwire sum_12_ ();
drwire sum_13_ ();
drwire sum_14_ ();
drwire sum_15_ ();
drwire sum_16_ ();
drwire sum_17_ ();
drwire sum_18_ ();
drwire sum_19_ ();
drwire sum_1_ ();
drwire sum_20_ ();
drwire sum_21_ ();
drwire sum_22_ ();
drwire sum_23_ ();
drwire sum_24_ ();
drwire sum_25_ ();
drwire sum_26_ ();
drwire sum_27_ ();
drwire sum_28_ ();
drwire sum_29_ ();
drwire sum_2_ ();
drwire sum_30_ ();
drwire sum_31_ ();
drwire sum_3_ ();
drwire sum_4_ ();
drwire sum_5_ ();
drwire sum_6_ ();
drwire sum_7_ ();
drwire sum_8_ ();
drwire sum_9_ ();
drwire v0_0_ ();
drwire v0_10_ ();
drwire v0_11_ ();
drwire v0_12_ ();
drwire v0_13_ ();
drwire v0_14_ ();
drwire v0_15_ ();
drwire v0_16_ ();
drwire v0_17_ ();
drwire v0_18_ ();
drwire v0_19_ ();
drwire v0_1_ ();
drwire v0_20_ ();
drwire v0_21_ ();
drwire v0_22_ ();
drwire v0_23_ ();
drwire v0_24_ ();
drwire v0_25_ ();
drwire v0_26_ ();
drwire v0_27_ ();
drwire v0_28_ ();
drwire v0_29_ ();
drwire v0_2_ ();
drwire v0_30_ ();
drwire v0_31_ ();
drwire v0_3_ ();
drwire v0_4_ ();
drwire v0_5_ ();
drwire v0_6_ ();
drwire v0_7_ ();
drwire v0_8_ ();
drwire v0_9_ ();
drwire v0_r_0_ ();
drwire v0_r_10_ ();
drwire v0_r_11_ ();
drwire v0_r_12_ ();
drwire v0_r_13_ ();
drwire v0_r_14_ ();
drwire v0_r_15_ ();
drwire v0_r_16_ ();
drwire v0_r_17_ ();
drwire v0_r_18_ ();
drwire v0_r_19_ ();
drwire v0_r_1_ ();
drwire v0_r_20_ ();
drwire v0_r_21_ ();
drwire v0_r_22_ ();
drwire v0_r_23_ ();
drwire v0_r_24_ ();
drwire v0_r_25_ ();
drwire v0_r_26_ ();
drwire v0_r_27_ ();
drwire v0_r_28_ ();
drwire v0_r_29_ ();
drwire v0_r_2_ ();
drwire v0_r_30_ ();
drwire v0_r_31_ ();
drwire v0_r_3_ ();
drwire v0_r_4_ ();
drwire v0_r_5_ ();
drwire v0_r_6_ ();
drwire v0_r_7_ ();
drwire v0_r_8_ ();
drwire v0_r_9_ ();
drwire v1_0_ ();
drwire v1_10_ ();
drwire v1_11_ ();
drwire v1_12_ ();
drwire v1_13_ ();
drwire v1_14_ ();
drwire v1_15_ ();
drwire v1_16_ ();
drwire v1_17_ ();
drwire v1_18_ ();
drwire v1_19_ ();
drwire v1_1_ ();
drwire v1_20_ ();
drwire v1_21_ ();
drwire v1_22_ ();
drwire v1_23_ ();
drwire v1_24_ ();
drwire v1_25_ ();
drwire v1_26_ ();
drwire v1_27_ ();
drwire v1_28_ ();
drwire v1_29_ ();
drwire v1_2_ ();
drwire v1_30_ ();
drwire v1_31_ ();
drwire v1_3_ ();
drwire v1_4_ ();
drwire v1_5_ ();
drwire v1_6_ ();
drwire v1_7_ ();
drwire v1_8_ ();
drwire v1_9_ ();
drwire v1_r_0_ ();
drwire v1_r_10_ ();
drwire v1_r_11_ ();
drwire v1_r_12_ ();
drwire v1_r_13_ ();
drwire v1_r_14_ ();
drwire v1_r_15_ ();
drwire v1_r_16_ ();
drwire v1_r_17_ ();
drwire v1_r_18_ ();
drwire v1_r_19_ ();
drwire v1_r_1_ ();
drwire v1_r_20_ ();
drwire v1_r_21_ ();
drwire v1_r_22_ ();
drwire v1_r_23_ ();
drwire v1_r_24_ ();
drwire v1_r_25_ ();
drwire v1_r_26_ ();
drwire v1_r_27_ ();
drwire v1_r_28_ ();
drwire v1_r_29_ ();
drwire v1_r_2_ ();
drwire v1_r_30_ ();
drwire v1_r_31_ ();
drwire v1_r_3_ ();
drwire v1_r_4_ ();
drwire v1_r_5_ ();
drwire v1_r_6_ ();
drwire v1_r_7_ ();
drwire v1_r_8_ ();
drwire v1_r_9_ ();
drwire in_enc_0 ();
drwire in_enc_1 ();
drwire in_enc_2 ();
drwire in_enc_3 ();
drwire in_enc_4 ();
drwire in_enc_5 ();
drwire in_enc_6 ();
drwire in_enc_7 ();
drwire in_enc_8 ();
drwire in_enc_9 ();
drwire in_enc_10 ();
drwire in_enc_11 ();
drwire in_enc_12 ();
drwire in_enc_13 ();
drwire in_enc_14 ();
drwire in_enc_15 ();
drwire in_enc_16 ();
drwire in_enc_17 ();
drwire in_enc_18 ();
drwire in_enc_19 ();
drwire in_enc_20 ();
drwire in_enc_21 ();
drwire in_enc_22 ();
drwire in_enc_23 ();
drwire in_enc_24 ();
drwire in_enc_25 ();
drwire in_enc_26 ();
drwire in_enc_27 ();
drwire in_enc_28 ();
drwire in_enc_29 ();
drwire in_enc_30 ();
drwire in_enc_31 ();
drwire in_enc_32 ();
drwire in_enc_33 ();
drwire in_enc_34 ();
drwire in_enc_35 ();
drwire in_enc_36 ();
drwire in_enc_37 ();
drwire in_enc_38 ();
drwire in_enc_39 ();
drwire in_enc_40 ();
drwire in_enc_41 ();
drwire in_enc_42 ();
drwire in_enc_43 ();
drwire in_enc_44 ();
drwire in_enc_45 ();
drwire in_enc_46 ();
drwire in_enc_47 ();
drwire in_enc_48 ();
drwire in_enc_49 ();
drwire in_enc_50 ();
drwire in_enc_51 ();
drwire in_enc_52 ();
drwire in_enc_53 ();
drwire in_enc_54 ();
drwire in_enc_55 ();
drwire in_enc_56 ();
drwire in_enc_57 ();
drwire in_enc_58 ();
drwire in_enc_59 ();
drwire in_enc_60 ();
drwire in_enc_61 ();
drwire in_enc_62 ();
drwire in_enc_63 ();
drwire out_enc_0 ();
drwire out_enc_1 ();
drwire out_enc_2 ();
drwire out_enc_3 ();
drwire out_enc_4 ();
drwire out_enc_5 ();
drwire out_enc_6 ();
drwire out_enc_7 ();
drwire out_enc_8 ();
drwire out_enc_9 ();
drwire out_enc_10 ();
drwire out_enc_11 ();
drwire out_enc_12 ();
drwire out_enc_13 ();
drwire out_enc_14 ();
drwire out_enc_15 ();
drwire out_enc_16 ();
drwire out_enc_17 ();
drwire out_enc_18 ();
drwire out_enc_19 ();
drwire out_enc_20 ();
drwire out_enc_21 ();
drwire out_enc_22 ();
drwire out_enc_23 ();
drwire out_enc_24 ();
drwire out_enc_25 ();
drwire out_enc_26 ();
drwire out_enc_27 ();
drwire out_enc_28 ();
drwire out_enc_29 ();
drwire out_enc_30 ();
drwire out_enc_31 ();
drwire out_enc_32 ();
drwire out_enc_33 ();
drwire out_enc_34 ();
drwire out_enc_35 ();
drwire out_enc_36 ();
drwire out_enc_37 ();
drwire out_enc_38 ();
drwire out_enc_39 ();
drwire out_enc_40 ();
drwire out_enc_41 ();
drwire out_enc_42 ();
drwire out_enc_43 ();
drwire out_enc_44 ();
drwire out_enc_45 ();
drwire out_enc_46 ();
drwire out_enc_47 ();
drwire out_enc_48 ();
drwire out_enc_49 ();
drwire out_enc_50 ();
drwire out_enc_51 ();
drwire out_enc_52 ();
drwire out_enc_53 ();
drwire out_enc_54 ();
drwire out_enc_55 ();
drwire out_enc_56 ();
drwire out_enc_57 ();
drwire out_enc_58 ();
drwire out_enc_59 ();
drwire out_enc_60 ();
drwire out_enc_61 ();
drwire out_enc_62 ();
drwire out_enc_63 ();
drwire key_0 ();
drwire key_1 ();
drwire key_2 ();
drwire key_3 ();
drwire key_4 ();
drwire key_5 ();
drwire key_6 ();
drwire key_7 ();
drwire key_8 ();
drwire key_9 ();
drwire key_10 ();
drwire key_11 ();
drwire key_12 ();
drwire key_13 ();
drwire key_14 ();
drwire key_15 ();
drwire key_16 ();
drwire key_17 ();
drwire key_18 ();
drwire key_19 ();
drwire key_20 ();
drwire key_21 ();
drwire key_22 ();
drwire key_23 ();
drwire key_24 ();
drwire key_25 ();
drwire key_26 ();
drwire key_27 ();
drwire key_28 ();
drwire key_29 ();
drwire key_30 ();
drwire key_31 ();
drwire key_32 ();
drwire key_33 ();
drwire key_34 ();
drwire key_35 ();
drwire key_36 ();
drwire key_37 ();
drwire key_38 ();
drwire key_39 ();
drwire key_40 ();
drwire key_41 ();
drwire key_42 ();
drwire key_43 ();
drwire key_44 ();
drwire key_45 ();
drwire key_46 ();
drwire key_47 ();
drwire key_48 ();
drwire key_49 ();
drwire key_50 ();
drwire key_51 ();
drwire key_52 ();
drwire key_53 ();
drwire key_54 ();
drwire key_55 ();
drwire key_56 ();
drwire key_57 ();
drwire key_58 ();
drwire key_59 ();
drwire key_60 ();
drwire key_61 ();
drwire key_62 ();
drwire key_63 ();
drwire key_64 ();
drwire key_65 ();
drwire key_66 ();
drwire key_67 ();
drwire key_68 ();
drwire key_69 ();
drwire key_70 ();
drwire key_71 ();
drwire key_72 ();
drwire key_73 ();
drwire key_74 ();
drwire key_75 ();
drwire key_76 ();
drwire key_77 ();
drwire key_78 ();
drwire key_79 ();
drwire key_80 ();
drwire key_81 ();
drwire key_82 ();
drwire key_83 ();
drwire key_84 ();
drwire key_85 ();
drwire key_86 ();
drwire key_87 ();
drwire key_88 ();
drwire key_89 ();
drwire key_90 ();
drwire key_91 ();
drwire key_92 ();
drwire key_93 ();
drwire key_94 ();
drwire key_95 ();
drwire key_96 ();
drwire key_97 ();
drwire key_98 ();
drwire key_99 ();
drwire key_100 ();
drwire key_101 ();
drwire key_102 ();
drwire key_103 ();
drwire key_104 ();
drwire key_105 ();
drwire key_106 ();
drwire key_107 ();
drwire key_108 ();
drwire key_109 ();
drwire key_110 ();
drwire key_111 ();
drwire key_112 ();
drwire key_113 ();
drwire key_114 ();
drwire key_115 ();
drwire key_116 ();
drwire key_117 ();
drwire key_118 ();
drwire key_119 ();
drwire key_120 ();
drwire key_121 ();
drwire key_122 ();
drwire key_123 ();
drwire key_124 ();
drwire key_125 ();
drwire key_126 ();
drwire key_127 ();
input  [63:0] in_enc_t, in_enc_f;
output [63:0] in_enc_ack;
drinput iin_enc_0 (.t(in_enc_t[0]), .f(in_enc_f[0]), .ack(in_enc_ack[0]), .drw(in_enc_0));
drinput iin_enc_1 (.t(in_enc_t[1]), .f(in_enc_f[1]), .ack(in_enc_ack[1]), .drw(in_enc_1));
drinput iin_enc_2 (.t(in_enc_t[2]), .f(in_enc_f[2]), .ack(in_enc_ack[2]), .drw(in_enc_2));
drinput iin_enc_3 (.t(in_enc_t[3]), .f(in_enc_f[3]), .ack(in_enc_ack[3]), .drw(in_enc_3));
drinput iin_enc_4 (.t(in_enc_t[4]), .f(in_enc_f[4]), .ack(in_enc_ack[4]), .drw(in_enc_4));
drinput iin_enc_5 (.t(in_enc_t[5]), .f(in_enc_f[5]), .ack(in_enc_ack[5]), .drw(in_enc_5));
drinput iin_enc_6 (.t(in_enc_t[6]), .f(in_enc_f[6]), .ack(in_enc_ack[6]), .drw(in_enc_6));
drinput iin_enc_7 (.t(in_enc_t[7]), .f(in_enc_f[7]), .ack(in_enc_ack[7]), .drw(in_enc_7));
drinput iin_enc_8 (.t(in_enc_t[8]), .f(in_enc_f[8]), .ack(in_enc_ack[8]), .drw(in_enc_8));
drinput iin_enc_9 (.t(in_enc_t[9]), .f(in_enc_f[9]), .ack(in_enc_ack[9]), .drw(in_enc_9));
drinput iin_enc_10 (.t(in_enc_t[10]), .f(in_enc_f[10]), .ack(in_enc_ack[10]), .drw(in_enc_10));
drinput iin_enc_11 (.t(in_enc_t[11]), .f(in_enc_f[11]), .ack(in_enc_ack[11]), .drw(in_enc_11));
drinput iin_enc_12 (.t(in_enc_t[12]), .f(in_enc_f[12]), .ack(in_enc_ack[12]), .drw(in_enc_12));
drinput iin_enc_13 (.t(in_enc_t[13]), .f(in_enc_f[13]), .ack(in_enc_ack[13]), .drw(in_enc_13));
drinput iin_enc_14 (.t(in_enc_t[14]), .f(in_enc_f[14]), .ack(in_enc_ack[14]), .drw(in_enc_14));
drinput iin_enc_15 (.t(in_enc_t[15]), .f(in_enc_f[15]), .ack(in_enc_ack[15]), .drw(in_enc_15));
drinput iin_enc_16 (.t(in_enc_t[16]), .f(in_enc_f[16]), .ack(in_enc_ack[16]), .drw(in_enc_16));
drinput iin_enc_17 (.t(in_enc_t[17]), .f(in_enc_f[17]), .ack(in_enc_ack[17]), .drw(in_enc_17));
drinput iin_enc_18 (.t(in_enc_t[18]), .f(in_enc_f[18]), .ack(in_enc_ack[18]), .drw(in_enc_18));
drinput iin_enc_19 (.t(in_enc_t[19]), .f(in_enc_f[19]), .ack(in_enc_ack[19]), .drw(in_enc_19));
drinput iin_enc_20 (.t(in_enc_t[20]), .f(in_enc_f[20]), .ack(in_enc_ack[20]), .drw(in_enc_20));
drinput iin_enc_21 (.t(in_enc_t[21]), .f(in_enc_f[21]), .ack(in_enc_ack[21]), .drw(in_enc_21));
drinput iin_enc_22 (.t(in_enc_t[22]), .f(in_enc_f[22]), .ack(in_enc_ack[22]), .drw(in_enc_22));
drinput iin_enc_23 (.t(in_enc_t[23]), .f(in_enc_f[23]), .ack(in_enc_ack[23]), .drw(in_enc_23));
drinput iin_enc_24 (.t(in_enc_t[24]), .f(in_enc_f[24]), .ack(in_enc_ack[24]), .drw(in_enc_24));
drinput iin_enc_25 (.t(in_enc_t[25]), .f(in_enc_f[25]), .ack(in_enc_ack[25]), .drw(in_enc_25));
drinput iin_enc_26 (.t(in_enc_t[26]), .f(in_enc_f[26]), .ack(in_enc_ack[26]), .drw(in_enc_26));
drinput iin_enc_27 (.t(in_enc_t[27]), .f(in_enc_f[27]), .ack(in_enc_ack[27]), .drw(in_enc_27));
drinput iin_enc_28 (.t(in_enc_t[28]), .f(in_enc_f[28]), .ack(in_enc_ack[28]), .drw(in_enc_28));
drinput iin_enc_29 (.t(in_enc_t[29]), .f(in_enc_f[29]), .ack(in_enc_ack[29]), .drw(in_enc_29));
drinput iin_enc_30 (.t(in_enc_t[30]), .f(in_enc_f[30]), .ack(in_enc_ack[30]), .drw(in_enc_30));
drinput iin_enc_31 (.t(in_enc_t[31]), .f(in_enc_f[31]), .ack(in_enc_ack[31]), .drw(in_enc_31));
drinput iin_enc_32 (.t(in_enc_t[32]), .f(in_enc_f[32]), .ack(in_enc_ack[32]), .drw(in_enc_32));
drinput iin_enc_33 (.t(in_enc_t[33]), .f(in_enc_f[33]), .ack(in_enc_ack[33]), .drw(in_enc_33));
drinput iin_enc_34 (.t(in_enc_t[34]), .f(in_enc_f[34]), .ack(in_enc_ack[34]), .drw(in_enc_34));
drinput iin_enc_35 (.t(in_enc_t[35]), .f(in_enc_f[35]), .ack(in_enc_ack[35]), .drw(in_enc_35));
drinput iin_enc_36 (.t(in_enc_t[36]), .f(in_enc_f[36]), .ack(in_enc_ack[36]), .drw(in_enc_36));
drinput iin_enc_37 (.t(in_enc_t[37]), .f(in_enc_f[37]), .ack(in_enc_ack[37]), .drw(in_enc_37));
drinput iin_enc_38 (.t(in_enc_t[38]), .f(in_enc_f[38]), .ack(in_enc_ack[38]), .drw(in_enc_38));
drinput iin_enc_39 (.t(in_enc_t[39]), .f(in_enc_f[39]), .ack(in_enc_ack[39]), .drw(in_enc_39));
drinput iin_enc_40 (.t(in_enc_t[40]), .f(in_enc_f[40]), .ack(in_enc_ack[40]), .drw(in_enc_40));
drinput iin_enc_41 (.t(in_enc_t[41]), .f(in_enc_f[41]), .ack(in_enc_ack[41]), .drw(in_enc_41));
drinput iin_enc_42 (.t(in_enc_t[42]), .f(in_enc_f[42]), .ack(in_enc_ack[42]), .drw(in_enc_42));
drinput iin_enc_43 (.t(in_enc_t[43]), .f(in_enc_f[43]), .ack(in_enc_ack[43]), .drw(in_enc_43));
drinput iin_enc_44 (.t(in_enc_t[44]), .f(in_enc_f[44]), .ack(in_enc_ack[44]), .drw(in_enc_44));
drinput iin_enc_45 (.t(in_enc_t[45]), .f(in_enc_f[45]), .ack(in_enc_ack[45]), .drw(in_enc_45));
drinput iin_enc_46 (.t(in_enc_t[46]), .f(in_enc_f[46]), .ack(in_enc_ack[46]), .drw(in_enc_46));
drinput iin_enc_47 (.t(in_enc_t[47]), .f(in_enc_f[47]), .ack(in_enc_ack[47]), .drw(in_enc_47));
drinput iin_enc_48 (.t(in_enc_t[48]), .f(in_enc_f[48]), .ack(in_enc_ack[48]), .drw(in_enc_48));
drinput iin_enc_49 (.t(in_enc_t[49]), .f(in_enc_f[49]), .ack(in_enc_ack[49]), .drw(in_enc_49));
drinput iin_enc_50 (.t(in_enc_t[50]), .f(in_enc_f[50]), .ack(in_enc_ack[50]), .drw(in_enc_50));
drinput iin_enc_51 (.t(in_enc_t[51]), .f(in_enc_f[51]), .ack(in_enc_ack[51]), .drw(in_enc_51));
drinput iin_enc_52 (.t(in_enc_t[52]), .f(in_enc_f[52]), .ack(in_enc_ack[52]), .drw(in_enc_52));
drinput iin_enc_53 (.t(in_enc_t[53]), .f(in_enc_f[53]), .ack(in_enc_ack[53]), .drw(in_enc_53));
drinput iin_enc_54 (.t(in_enc_t[54]), .f(in_enc_f[54]), .ack(in_enc_ack[54]), .drw(in_enc_54));
drinput iin_enc_55 (.t(in_enc_t[55]), .f(in_enc_f[55]), .ack(in_enc_ack[55]), .drw(in_enc_55));
drinput iin_enc_56 (.t(in_enc_t[56]), .f(in_enc_f[56]), .ack(in_enc_ack[56]), .drw(in_enc_56));
drinput iin_enc_57 (.t(in_enc_t[57]), .f(in_enc_f[57]), .ack(in_enc_ack[57]), .drw(in_enc_57));
drinput iin_enc_58 (.t(in_enc_t[58]), .f(in_enc_f[58]), .ack(in_enc_ack[58]), .drw(in_enc_58));
drinput iin_enc_59 (.t(in_enc_t[59]), .f(in_enc_f[59]), .ack(in_enc_ack[59]), .drw(in_enc_59));
drinput iin_enc_60 (.t(in_enc_t[60]), .f(in_enc_f[60]), .ack(in_enc_ack[60]), .drw(in_enc_60));
drinput iin_enc_61 (.t(in_enc_t[61]), .f(in_enc_f[61]), .ack(in_enc_ack[61]), .drw(in_enc_61));
drinput iin_enc_62 (.t(in_enc_t[62]), .f(in_enc_f[62]), .ack(in_enc_ack[62]), .drw(in_enc_62));
drinput iin_enc_63 (.t(in_enc_t[63]), .f(in_enc_f[63]), .ack(in_enc_ack[63]), .drw(in_enc_63));
input  [127:0] key_t, key_f;
output [127:0] key_ack;
drinput ikey_0 (.t(key_t[0]), .f(key_f[0]), .ack(key_ack[0]), .drw(key_0));
drinput ikey_1 (.t(key_t[1]), .f(key_f[1]), .ack(key_ack[1]), .drw(key_1));
drinput ikey_2 (.t(key_t[2]), .f(key_f[2]), .ack(key_ack[2]), .drw(key_2));
drinput ikey_3 (.t(key_t[3]), .f(key_f[3]), .ack(key_ack[3]), .drw(key_3));
drinput ikey_4 (.t(key_t[4]), .f(key_f[4]), .ack(key_ack[4]), .drw(key_4));
drinput ikey_5 (.t(key_t[5]), .f(key_f[5]), .ack(key_ack[5]), .drw(key_5));
drinput ikey_6 (.t(key_t[6]), .f(key_f[6]), .ack(key_ack[6]), .drw(key_6));
drinput ikey_7 (.t(key_t[7]), .f(key_f[7]), .ack(key_ack[7]), .drw(key_7));
drinput ikey_8 (.t(key_t[8]), .f(key_f[8]), .ack(key_ack[8]), .drw(key_8));
drinput ikey_9 (.t(key_t[9]), .f(key_f[9]), .ack(key_ack[9]), .drw(key_9));
drinput ikey_10 (.t(key_t[10]), .f(key_f[10]), .ack(key_ack[10]), .drw(key_10));
drinput ikey_11 (.t(key_t[11]), .f(key_f[11]), .ack(key_ack[11]), .drw(key_11));
drinput ikey_12 (.t(key_t[12]), .f(key_f[12]), .ack(key_ack[12]), .drw(key_12));
drinput ikey_13 (.t(key_t[13]), .f(key_f[13]), .ack(key_ack[13]), .drw(key_13));
drinput ikey_14 (.t(key_t[14]), .f(key_f[14]), .ack(key_ack[14]), .drw(key_14));
drinput ikey_15 (.t(key_t[15]), .f(key_f[15]), .ack(key_ack[15]), .drw(key_15));
drinput ikey_16 (.t(key_t[16]), .f(key_f[16]), .ack(key_ack[16]), .drw(key_16));
drinput ikey_17 (.t(key_t[17]), .f(key_f[17]), .ack(key_ack[17]), .drw(key_17));
drinput ikey_18 (.t(key_t[18]), .f(key_f[18]), .ack(key_ack[18]), .drw(key_18));
drinput ikey_19 (.t(key_t[19]), .f(key_f[19]), .ack(key_ack[19]), .drw(key_19));
drinput ikey_20 (.t(key_t[20]), .f(key_f[20]), .ack(key_ack[20]), .drw(key_20));
drinput ikey_21 (.t(key_t[21]), .f(key_f[21]), .ack(key_ack[21]), .drw(key_21));
drinput ikey_22 (.t(key_t[22]), .f(key_f[22]), .ack(key_ack[22]), .drw(key_22));
drinput ikey_23 (.t(key_t[23]), .f(key_f[23]), .ack(key_ack[23]), .drw(key_23));
drinput ikey_24 (.t(key_t[24]), .f(key_f[24]), .ack(key_ack[24]), .drw(key_24));
drinput ikey_25 (.t(key_t[25]), .f(key_f[25]), .ack(key_ack[25]), .drw(key_25));
drinput ikey_26 (.t(key_t[26]), .f(key_f[26]), .ack(key_ack[26]), .drw(key_26));
drinput ikey_27 (.t(key_t[27]), .f(key_f[27]), .ack(key_ack[27]), .drw(key_27));
drinput ikey_28 (.t(key_t[28]), .f(key_f[28]), .ack(key_ack[28]), .drw(key_28));
drinput ikey_29 (.t(key_t[29]), .f(key_f[29]), .ack(key_ack[29]), .drw(key_29));
drinput ikey_30 (.t(key_t[30]), .f(key_f[30]), .ack(key_ack[30]), .drw(key_30));
drinput ikey_31 (.t(key_t[31]), .f(key_f[31]), .ack(key_ack[31]), .drw(key_31));
drinput ikey_32 (.t(key_t[32]), .f(key_f[32]), .ack(key_ack[32]), .drw(key_32));
drinput ikey_33 (.t(key_t[33]), .f(key_f[33]), .ack(key_ack[33]), .drw(key_33));
drinput ikey_34 (.t(key_t[34]), .f(key_f[34]), .ack(key_ack[34]), .drw(key_34));
drinput ikey_35 (.t(key_t[35]), .f(key_f[35]), .ack(key_ack[35]), .drw(key_35));
drinput ikey_36 (.t(key_t[36]), .f(key_f[36]), .ack(key_ack[36]), .drw(key_36));
drinput ikey_37 (.t(key_t[37]), .f(key_f[37]), .ack(key_ack[37]), .drw(key_37));
drinput ikey_38 (.t(key_t[38]), .f(key_f[38]), .ack(key_ack[38]), .drw(key_38));
drinput ikey_39 (.t(key_t[39]), .f(key_f[39]), .ack(key_ack[39]), .drw(key_39));
drinput ikey_40 (.t(key_t[40]), .f(key_f[40]), .ack(key_ack[40]), .drw(key_40));
drinput ikey_41 (.t(key_t[41]), .f(key_f[41]), .ack(key_ack[41]), .drw(key_41));
drinput ikey_42 (.t(key_t[42]), .f(key_f[42]), .ack(key_ack[42]), .drw(key_42));
drinput ikey_43 (.t(key_t[43]), .f(key_f[43]), .ack(key_ack[43]), .drw(key_43));
drinput ikey_44 (.t(key_t[44]), .f(key_f[44]), .ack(key_ack[44]), .drw(key_44));
drinput ikey_45 (.t(key_t[45]), .f(key_f[45]), .ack(key_ack[45]), .drw(key_45));
drinput ikey_46 (.t(key_t[46]), .f(key_f[46]), .ack(key_ack[46]), .drw(key_46));
drinput ikey_47 (.t(key_t[47]), .f(key_f[47]), .ack(key_ack[47]), .drw(key_47));
drinput ikey_48 (.t(key_t[48]), .f(key_f[48]), .ack(key_ack[48]), .drw(key_48));
drinput ikey_49 (.t(key_t[49]), .f(key_f[49]), .ack(key_ack[49]), .drw(key_49));
drinput ikey_50 (.t(key_t[50]), .f(key_f[50]), .ack(key_ack[50]), .drw(key_50));
drinput ikey_51 (.t(key_t[51]), .f(key_f[51]), .ack(key_ack[51]), .drw(key_51));
drinput ikey_52 (.t(key_t[52]), .f(key_f[52]), .ack(key_ack[52]), .drw(key_52));
drinput ikey_53 (.t(key_t[53]), .f(key_f[53]), .ack(key_ack[53]), .drw(key_53));
drinput ikey_54 (.t(key_t[54]), .f(key_f[54]), .ack(key_ack[54]), .drw(key_54));
drinput ikey_55 (.t(key_t[55]), .f(key_f[55]), .ack(key_ack[55]), .drw(key_55));
drinput ikey_56 (.t(key_t[56]), .f(key_f[56]), .ack(key_ack[56]), .drw(key_56));
drinput ikey_57 (.t(key_t[57]), .f(key_f[57]), .ack(key_ack[57]), .drw(key_57));
drinput ikey_58 (.t(key_t[58]), .f(key_f[58]), .ack(key_ack[58]), .drw(key_58));
drinput ikey_59 (.t(key_t[59]), .f(key_f[59]), .ack(key_ack[59]), .drw(key_59));
drinput ikey_60 (.t(key_t[60]), .f(key_f[60]), .ack(key_ack[60]), .drw(key_60));
drinput ikey_61 (.t(key_t[61]), .f(key_f[61]), .ack(key_ack[61]), .drw(key_61));
drinput ikey_62 (.t(key_t[62]), .f(key_f[62]), .ack(key_ack[62]), .drw(key_62));
drinput ikey_63 (.t(key_t[63]), .f(key_f[63]), .ack(key_ack[63]), .drw(key_63));
drinput ikey_64 (.t(key_t[64]), .f(key_f[64]), .ack(key_ack[64]), .drw(key_64));
drinput ikey_65 (.t(key_t[65]), .f(key_f[65]), .ack(key_ack[65]), .drw(key_65));
drinput ikey_66 (.t(key_t[66]), .f(key_f[66]), .ack(key_ack[66]), .drw(key_66));
drinput ikey_67 (.t(key_t[67]), .f(key_f[67]), .ack(key_ack[67]), .drw(key_67));
drinput ikey_68 (.t(key_t[68]), .f(key_f[68]), .ack(key_ack[68]), .drw(key_68));
drinput ikey_69 (.t(key_t[69]), .f(key_f[69]), .ack(key_ack[69]), .drw(key_69));
drinput ikey_70 (.t(key_t[70]), .f(key_f[70]), .ack(key_ack[70]), .drw(key_70));
drinput ikey_71 (.t(key_t[71]), .f(key_f[71]), .ack(key_ack[71]), .drw(key_71));
drinput ikey_72 (.t(key_t[72]), .f(key_f[72]), .ack(key_ack[72]), .drw(key_72));
drinput ikey_73 (.t(key_t[73]), .f(key_f[73]), .ack(key_ack[73]), .drw(key_73));
drinput ikey_74 (.t(key_t[74]), .f(key_f[74]), .ack(key_ack[74]), .drw(key_74));
drinput ikey_75 (.t(key_t[75]), .f(key_f[75]), .ack(key_ack[75]), .drw(key_75));
drinput ikey_76 (.t(key_t[76]), .f(key_f[76]), .ack(key_ack[76]), .drw(key_76));
drinput ikey_77 (.t(key_t[77]), .f(key_f[77]), .ack(key_ack[77]), .drw(key_77));
drinput ikey_78 (.t(key_t[78]), .f(key_f[78]), .ack(key_ack[78]), .drw(key_78));
drinput ikey_79 (.t(key_t[79]), .f(key_f[79]), .ack(key_ack[79]), .drw(key_79));
drinput ikey_80 (.t(key_t[80]), .f(key_f[80]), .ack(key_ack[80]), .drw(key_80));
drinput ikey_81 (.t(key_t[81]), .f(key_f[81]), .ack(key_ack[81]), .drw(key_81));
drinput ikey_82 (.t(key_t[82]), .f(key_f[82]), .ack(key_ack[82]), .drw(key_82));
drinput ikey_83 (.t(key_t[83]), .f(key_f[83]), .ack(key_ack[83]), .drw(key_83));
drinput ikey_84 (.t(key_t[84]), .f(key_f[84]), .ack(key_ack[84]), .drw(key_84));
drinput ikey_85 (.t(key_t[85]), .f(key_f[85]), .ack(key_ack[85]), .drw(key_85));
drinput ikey_86 (.t(key_t[86]), .f(key_f[86]), .ack(key_ack[86]), .drw(key_86));
drinput ikey_87 (.t(key_t[87]), .f(key_f[87]), .ack(key_ack[87]), .drw(key_87));
drinput ikey_88 (.t(key_t[88]), .f(key_f[88]), .ack(key_ack[88]), .drw(key_88));
drinput ikey_89 (.t(key_t[89]), .f(key_f[89]), .ack(key_ack[89]), .drw(key_89));
drinput ikey_90 (.t(key_t[90]), .f(key_f[90]), .ack(key_ack[90]), .drw(key_90));
drinput ikey_91 (.t(key_t[91]), .f(key_f[91]), .ack(key_ack[91]), .drw(key_91));
drinput ikey_92 (.t(key_t[92]), .f(key_f[92]), .ack(key_ack[92]), .drw(key_92));
drinput ikey_93 (.t(key_t[93]), .f(key_f[93]), .ack(key_ack[93]), .drw(key_93));
drinput ikey_94 (.t(key_t[94]), .f(key_f[94]), .ack(key_ack[94]), .drw(key_94));
drinput ikey_95 (.t(key_t[95]), .f(key_f[95]), .ack(key_ack[95]), .drw(key_95));
drinput ikey_96 (.t(key_t[96]), .f(key_f[96]), .ack(key_ack[96]), .drw(key_96));
drinput ikey_97 (.t(key_t[97]), .f(key_f[97]), .ack(key_ack[97]), .drw(key_97));
drinput ikey_98 (.t(key_t[98]), .f(key_f[98]), .ack(key_ack[98]), .drw(key_98));
drinput ikey_99 (.t(key_t[99]), .f(key_f[99]), .ack(key_ack[99]), .drw(key_99));
drinput ikey_100 (.t(key_t[100]), .f(key_f[100]), .ack(key_ack[100]), .drw(key_100));
drinput ikey_101 (.t(key_t[101]), .f(key_f[101]), .ack(key_ack[101]), .drw(key_101));
drinput ikey_102 (.t(key_t[102]), .f(key_f[102]), .ack(key_ack[102]), .drw(key_102));
drinput ikey_103 (.t(key_t[103]), .f(key_f[103]), .ack(key_ack[103]), .drw(key_103));
drinput ikey_104 (.t(key_t[104]), .f(key_f[104]), .ack(key_ack[104]), .drw(key_104));
drinput ikey_105 (.t(key_t[105]), .f(key_f[105]), .ack(key_ack[105]), .drw(key_105));
drinput ikey_106 (.t(key_t[106]), .f(key_f[106]), .ack(key_ack[106]), .drw(key_106));
drinput ikey_107 (.t(key_t[107]), .f(key_f[107]), .ack(key_ack[107]), .drw(key_107));
drinput ikey_108 (.t(key_t[108]), .f(key_f[108]), .ack(key_ack[108]), .drw(key_108));
drinput ikey_109 (.t(key_t[109]), .f(key_f[109]), .ack(key_ack[109]), .drw(key_109));
drinput ikey_110 (.t(key_t[110]), .f(key_f[110]), .ack(key_ack[110]), .drw(key_110));
drinput ikey_111 (.t(key_t[111]), .f(key_f[111]), .ack(key_ack[111]), .drw(key_111));
drinput ikey_112 (.t(key_t[112]), .f(key_f[112]), .ack(key_ack[112]), .drw(key_112));
drinput ikey_113 (.t(key_t[113]), .f(key_f[113]), .ack(key_ack[113]), .drw(key_113));
drinput ikey_114 (.t(key_t[114]), .f(key_f[114]), .ack(key_ack[114]), .drw(key_114));
drinput ikey_115 (.t(key_t[115]), .f(key_f[115]), .ack(key_ack[115]), .drw(key_115));
drinput ikey_116 (.t(key_t[116]), .f(key_f[116]), .ack(key_ack[116]), .drw(key_116));
drinput ikey_117 (.t(key_t[117]), .f(key_f[117]), .ack(key_ack[117]), .drw(key_117));
drinput ikey_118 (.t(key_t[118]), .f(key_f[118]), .ack(key_ack[118]), .drw(key_118));
drinput ikey_119 (.t(key_t[119]), .f(key_f[119]), .ack(key_ack[119]), .drw(key_119));
drinput ikey_120 (.t(key_t[120]), .f(key_f[120]), .ack(key_ack[120]), .drw(key_120));
drinput ikey_121 (.t(key_t[121]), .f(key_f[121]), .ack(key_ack[121]), .drw(key_121));
drinput ikey_122 (.t(key_t[122]), .f(key_f[122]), .ack(key_ack[122]), .drw(key_122));
drinput ikey_123 (.t(key_t[123]), .f(key_f[123]), .ack(key_ack[123]), .drw(key_123));
drinput ikey_124 (.t(key_t[124]), .f(key_f[124]), .ack(key_ack[124]), .drw(key_124));
drinput ikey_125 (.t(key_t[125]), .f(key_f[125]), .ack(key_ack[125]), .drw(key_125));
drinput ikey_126 (.t(key_t[126]), .f(key_f[126]), .ack(key_ack[126]), .drw(key_126));
drinput ikey_127 (.t(key_t[127]), .f(key_f[127]), .ack(key_ack[127]), .drw(key_127));
output [63:0] out_enc_t, out_enc_f;
input  [63:0] out_enc_ack;
droutput iout_enc_0 (.t(out_enc_t[0]), .f(out_enc_f[0]), .ack(out_enc_ack[0]), .drw(out_enc_0));
droutput iout_enc_1 (.t(out_enc_t[1]), .f(out_enc_f[1]), .ack(out_enc_ack[1]), .drw(out_enc_1));
droutput iout_enc_2 (.t(out_enc_t[2]), .f(out_enc_f[2]), .ack(out_enc_ack[2]), .drw(out_enc_2));
droutput iout_enc_3 (.t(out_enc_t[3]), .f(out_enc_f[3]), .ack(out_enc_ack[3]), .drw(out_enc_3));
droutput iout_enc_4 (.t(out_enc_t[4]), .f(out_enc_f[4]), .ack(out_enc_ack[4]), .drw(out_enc_4));
droutput iout_enc_5 (.t(out_enc_t[5]), .f(out_enc_f[5]), .ack(out_enc_ack[5]), .drw(out_enc_5));
droutput iout_enc_6 (.t(out_enc_t[6]), .f(out_enc_f[6]), .ack(out_enc_ack[6]), .drw(out_enc_6));
droutput iout_enc_7 (.t(out_enc_t[7]), .f(out_enc_f[7]), .ack(out_enc_ack[7]), .drw(out_enc_7));
droutput iout_enc_8 (.t(out_enc_t[8]), .f(out_enc_f[8]), .ack(out_enc_ack[8]), .drw(out_enc_8));
droutput iout_enc_9 (.t(out_enc_t[9]), .f(out_enc_f[9]), .ack(out_enc_ack[9]), .drw(out_enc_9));
droutput iout_enc_10 (.t(out_enc_t[10]), .f(out_enc_f[10]), .ack(out_enc_ack[10]), .drw(out_enc_10));
droutput iout_enc_11 (.t(out_enc_t[11]), .f(out_enc_f[11]), .ack(out_enc_ack[11]), .drw(out_enc_11));
droutput iout_enc_12 (.t(out_enc_t[12]), .f(out_enc_f[12]), .ack(out_enc_ack[12]), .drw(out_enc_12));
droutput iout_enc_13 (.t(out_enc_t[13]), .f(out_enc_f[13]), .ack(out_enc_ack[13]), .drw(out_enc_13));
droutput iout_enc_14 (.t(out_enc_t[14]), .f(out_enc_f[14]), .ack(out_enc_ack[14]), .drw(out_enc_14));
droutput iout_enc_15 (.t(out_enc_t[15]), .f(out_enc_f[15]), .ack(out_enc_ack[15]), .drw(out_enc_15));
droutput iout_enc_16 (.t(out_enc_t[16]), .f(out_enc_f[16]), .ack(out_enc_ack[16]), .drw(out_enc_16));
droutput iout_enc_17 (.t(out_enc_t[17]), .f(out_enc_f[17]), .ack(out_enc_ack[17]), .drw(out_enc_17));
droutput iout_enc_18 (.t(out_enc_t[18]), .f(out_enc_f[18]), .ack(out_enc_ack[18]), .drw(out_enc_18));
droutput iout_enc_19 (.t(out_enc_t[19]), .f(out_enc_f[19]), .ack(out_enc_ack[19]), .drw(out_enc_19));
droutput iout_enc_20 (.t(out_enc_t[20]), .f(out_enc_f[20]), .ack(out_enc_ack[20]), .drw(out_enc_20));
droutput iout_enc_21 (.t(out_enc_t[21]), .f(out_enc_f[21]), .ack(out_enc_ack[21]), .drw(out_enc_21));
droutput iout_enc_22 (.t(out_enc_t[22]), .f(out_enc_f[22]), .ack(out_enc_ack[22]), .drw(out_enc_22));
droutput iout_enc_23 (.t(out_enc_t[23]), .f(out_enc_f[23]), .ack(out_enc_ack[23]), .drw(out_enc_23));
droutput iout_enc_24 (.t(out_enc_t[24]), .f(out_enc_f[24]), .ack(out_enc_ack[24]), .drw(out_enc_24));
droutput iout_enc_25 (.t(out_enc_t[25]), .f(out_enc_f[25]), .ack(out_enc_ack[25]), .drw(out_enc_25));
droutput iout_enc_26 (.t(out_enc_t[26]), .f(out_enc_f[26]), .ack(out_enc_ack[26]), .drw(out_enc_26));
droutput iout_enc_27 (.t(out_enc_t[27]), .f(out_enc_f[27]), .ack(out_enc_ack[27]), .drw(out_enc_27));
droutput iout_enc_28 (.t(out_enc_t[28]), .f(out_enc_f[28]), .ack(out_enc_ack[28]), .drw(out_enc_28));
droutput iout_enc_29 (.t(out_enc_t[29]), .f(out_enc_f[29]), .ack(out_enc_ack[29]), .drw(out_enc_29));
droutput iout_enc_30 (.t(out_enc_t[30]), .f(out_enc_f[30]), .ack(out_enc_ack[30]), .drw(out_enc_30));
droutput iout_enc_31 (.t(out_enc_t[31]), .f(out_enc_f[31]), .ack(out_enc_ack[31]), .drw(out_enc_31));
droutput iout_enc_32 (.t(out_enc_t[32]), .f(out_enc_f[32]), .ack(out_enc_ack[32]), .drw(out_enc_32));
droutput iout_enc_33 (.t(out_enc_t[33]), .f(out_enc_f[33]), .ack(out_enc_ack[33]), .drw(out_enc_33));
droutput iout_enc_34 (.t(out_enc_t[34]), .f(out_enc_f[34]), .ack(out_enc_ack[34]), .drw(out_enc_34));
droutput iout_enc_35 (.t(out_enc_t[35]), .f(out_enc_f[35]), .ack(out_enc_ack[35]), .drw(out_enc_35));
droutput iout_enc_36 (.t(out_enc_t[36]), .f(out_enc_f[36]), .ack(out_enc_ack[36]), .drw(out_enc_36));
droutput iout_enc_37 (.t(out_enc_t[37]), .f(out_enc_f[37]), .ack(out_enc_ack[37]), .drw(out_enc_37));
droutput iout_enc_38 (.t(out_enc_t[38]), .f(out_enc_f[38]), .ack(out_enc_ack[38]), .drw(out_enc_38));
droutput iout_enc_39 (.t(out_enc_t[39]), .f(out_enc_f[39]), .ack(out_enc_ack[39]), .drw(out_enc_39));
droutput iout_enc_40 (.t(out_enc_t[40]), .f(out_enc_f[40]), .ack(out_enc_ack[40]), .drw(out_enc_40));
droutput iout_enc_41 (.t(out_enc_t[41]), .f(out_enc_f[41]), .ack(out_enc_ack[41]), .drw(out_enc_41));
droutput iout_enc_42 (.t(out_enc_t[42]), .f(out_enc_f[42]), .ack(out_enc_ack[42]), .drw(out_enc_42));
droutput iout_enc_43 (.t(out_enc_t[43]), .f(out_enc_f[43]), .ack(out_enc_ack[43]), .drw(out_enc_43));
droutput iout_enc_44 (.t(out_enc_t[44]), .f(out_enc_f[44]), .ack(out_enc_ack[44]), .drw(out_enc_44));
droutput iout_enc_45 (.t(out_enc_t[45]), .f(out_enc_f[45]), .ack(out_enc_ack[45]), .drw(out_enc_45));
droutput iout_enc_46 (.t(out_enc_t[46]), .f(out_enc_f[46]), .ack(out_enc_ack[46]), .drw(out_enc_46));
droutput iout_enc_47 (.t(out_enc_t[47]), .f(out_enc_f[47]), .ack(out_enc_ack[47]), .drw(out_enc_47));
droutput iout_enc_48 (.t(out_enc_t[48]), .f(out_enc_f[48]), .ack(out_enc_ack[48]), .drw(out_enc_48));
droutput iout_enc_49 (.t(out_enc_t[49]), .f(out_enc_f[49]), .ack(out_enc_ack[49]), .drw(out_enc_49));
droutput iout_enc_50 (.t(out_enc_t[50]), .f(out_enc_f[50]), .ack(out_enc_ack[50]), .drw(out_enc_50));
droutput iout_enc_51 (.t(out_enc_t[51]), .f(out_enc_f[51]), .ack(out_enc_ack[51]), .drw(out_enc_51));
droutput iout_enc_52 (.t(out_enc_t[52]), .f(out_enc_f[52]), .ack(out_enc_ack[52]), .drw(out_enc_52));
droutput iout_enc_53 (.t(out_enc_t[53]), .f(out_enc_f[53]), .ack(out_enc_ack[53]), .drw(out_enc_53));
droutput iout_enc_54 (.t(out_enc_t[54]), .f(out_enc_f[54]), .ack(out_enc_ack[54]), .drw(out_enc_54));
droutput iout_enc_55 (.t(out_enc_t[55]), .f(out_enc_f[55]), .ack(out_enc_ack[55]), .drw(out_enc_55));
droutput iout_enc_56 (.t(out_enc_t[56]), .f(out_enc_f[56]), .ack(out_enc_ack[56]), .drw(out_enc_56));
droutput iout_enc_57 (.t(out_enc_t[57]), .f(out_enc_f[57]), .ack(out_enc_ack[57]), .drw(out_enc_57));
droutput iout_enc_58 (.t(out_enc_t[58]), .f(out_enc_f[58]), .ack(out_enc_ack[58]), .drw(out_enc_58));
droutput iout_enc_59 (.t(out_enc_t[59]), .f(out_enc_f[59]), .ack(out_enc_ack[59]), .drw(out_enc_59));
droutput iout_enc_60 (.t(out_enc_t[60]), .f(out_enc_f[60]), .ack(out_enc_ack[60]), .drw(out_enc_60));
droutput iout_enc_61 (.t(out_enc_t[61]), .f(out_enc_f[61]), .ack(out_enc_ack[61]), .drw(out_enc_61));
droutput iout_enc_62 (.t(out_enc_t[62]), .f(out_enc_f[62]), .ack(out_enc_ack[62]), .drw(out_enc_62));
droutput iout_enc_63 (.t(out_enc_t[63]), .f(out_enc_f[63]), .ack(out_enc_ack[63]), .drw(out_enc_63));
xor2 g2841__8780 (.a(n_2033), .b(n_1998), .y(n_974));
xor2 g2844__1474 (.a(n_3490), .b(n_1239), .y(n_981));
xor2 g2846__9682 (.a(n_1216), .b(n_3505), .y(n_967));
xor2 g2847__2683 (.a(n_1998), .b(n_1241), .y(n_983));
xor2 g2850__2900 (.a(n_1224), .b(n_3708), .y(n_975));
xor2 g2851__2391 (.a(n_3580), .b(n_1243), .y(n_985));
xor2 g2854__8757 (.a(n_2005), .b(n_1245), .y(n_987));
xor2 g2855__1786 (.a(n_2961), .b(n_1246), .y(n_988));
xor2 g2856__5953 (.a(n_1217), .b(n_4306), .y(n_968));
xor2 g2858__7114 (.a(n_1235), .b(n_1244), .y(n_986));
zbuf g361__7344 (.a(v0_6_), .en(n_645), .y(out_enc_38));
zbuf g346__1840 (.a(v0_26_), .en(n_645), .y(out_enc_58));
zbuf g347__5019 (.a(v0_25_), .en(n_645), .y(out_enc_57));
zbuf g357__1857 (.a(v0_10_), .en(n_645), .y(out_enc_42));
zbuf g358__9906 (.a(v0_9_), .en(n_645), .y(out_enc_41));
zbuf g389__8780 (.a(v1_10_), .en(n_645), .y(out_enc_10));
zbuf g390__4296 (.a(v1_9_), .en(n_645), .y(out_enc_9));
zbuf g391__3772 (.a(v1_8_), .en(n_645), .y(out_enc_8));
zbuf g392__1474 (.a(v1_7_), .en(n_645), .y(out_enc_7));
zbuf g359__4547 (.a(v0_8_), .en(n_645), .y(out_enc_40));
zbuf g393__9682 (.a(v1_6_), .en(n_645), .y(out_enc_6));
zbuf g394__2683 (.a(v1_5_), .en(n_645), .y(out_enc_5));
zbuf g360__1309 (.a(v0_7_), .en(n_645), .y(out_enc_39));
zbuf g395__6877 (.a(v1_4_), .en(n_645), .y(out_enc_4));
zbuf g396__2900 (.a(v1_3_), .en(n_645), .y(out_enc_3));
zbuf g348__2391 (.a(v0_24_), .en(n_645), .y(out_enc_56));
zbuf g341__7675 (.a(v0_31_), .en(n_645), .y(out_enc_63));
zbuf g397__7118 (.a(v1_2_), .en(n_645), .y(out_enc_2));
zbuf g398__8757 (.a(v1_1_), .en(n_645), .y(out_enc_1));
zbuf g362__1786 (.a(v0_5_), .en(n_645), .y(out_enc_37));
zbuf g399__5953 (.a(v1_0_), .en(n_645), .y(out_enc_0));
zbuf g349__5703 (.a(v0_23_), .en(n_645), .y(out_enc_55));
zbuf g363__7114 (.a(v0_4_), .en(n_645), .y(out_enc_36));
zbuf g364__5266 (.a(v0_3_), .en(n_645), .y(out_enc_35));
zbuf g350__2250 (.a(v0_22_), .en(n_645), .y(out_enc_54));
zbuf g11__6083 (.a(v0_21_), .en(n_645), .y(out_enc_53));
zbuf g365__2703 (.a(v0_2_), .en(n_645), .y(out_enc_34));
zbuf g366__5795 (.a(v0_1_), .en(n_645), .y(out_enc_33));
zbuf g367__7344 (.a(v0_0_), .en(n_645), .y(out_enc_32));
zbuf g368__1840 (.a(v1_31_), .en(n_645), .y(out_enc_31));
zbuf g12__5019 (.a(v0_20_), .en(n_645), .y(out_enc_52));
zbuf g369__1857 (.a(v1_30_), .en(n_645), .y(out_enc_30));
zbuf g379__9906 (.a(v1_20_), .en(n_645), .y(out_enc_20));
zbuf g13__8780 (.a(v0_19_), .en(n_645), .y(out_enc_51));
zbuf g371__4296 (.a(v1_28_), .en(n_645), .y(out_enc_28));
zbuf g372__3772 (.a(v1_27_), .en(n_645), .y(out_enc_27));
zbuf g342__1474 (.a(v0_30_), .en(n_645), .y(out_enc_62));
zbuf g343__4547 (.a(v0_29_), .en(n_645), .y(out_enc_61));
zbuf g14__9682 (.a(v0_18_), .en(n_645), .y(out_enc_50));
zbuf g373__2683 (.a(v1_26_), .en(n_645), .y(out_enc_26));
zbuf g374__1309 (.a(v1_25_), .en(n_645), .y(out_enc_25));
zbuf g15__6877 (.a(v0_17_), .en(n_645), .y(out_enc_49));
zbuf g375__2900 (.a(v1_24_), .en(n_645), .y(out_enc_24));
zbuf g376__2391 (.a(v1_23_), .en(n_645), .y(out_enc_23));
zbuf g351__7675 (.a(v0_16_), .en(n_645), .y(out_enc_48));
zbuf g377__7118 (.a(v1_22_), .en(n_645), .y(out_enc_22));
zbuf g378__8757 (.a(v1_21_), .en(n_645), .y(out_enc_21));
zbuf g352__1786 (.a(v0_15_), .en(n_645), .y(out_enc_47));
zbuf g370__5953 (.a(v1_29_), .en(n_645), .y(out_enc_29));
zbuf g380__5703 (.a(v1_19_), .en(n_645), .y(out_enc_19));
zbuf g344__7114 (.a(v0_28_), .en(n_645), .y(out_enc_60));
zbuf g353__5266 (.a(v0_14_), .en(n_645), .y(out_enc_46));
zbuf g381__2250 (.a(v1_18_), .en(n_645), .y(out_enc_18));
zbuf g382__6083 (.a(v1_17_), .en(n_645), .y(out_enc_17));
zbuf g354__2703 (.a(v0_13_), .en(n_645), .y(out_enc_45));
zbuf g383__5795 (.a(v1_16_), .en(n_645), .y(out_enc_16));
zbuf g384__7344 (.a(v1_15_), .en(n_645), .y(out_enc_15));
zbuf g345__1840 (.a(v0_27_), .en(n_645), .y(out_enc_59));
zbuf g355__5019 (.a(v0_12_), .en(n_645), .y(out_enc_44));
zbuf g385__1857 (.a(v1_14_), .en(n_645), .y(out_enc_14));
zbuf g386__9906 (.a(v1_13_), .en(n_645), .y(out_enc_13));
zbuf g356__8780 (.a(v0_11_), .en(n_645), .y(out_enc_43));
zbuf g387__4296 (.a(v1_12_), .en(n_645), .y(out_enc_12));
zbuf g388__3772 (.a(v1_11_), .en(n_645), .y(out_enc_11));
inv g5820 (.a(n_645), .y(n_647));
nor2 g5821__1474 (.a(n_649), .b(counter_10_), .y(n_645));
inv g5822 (.a(n_644), .y(n_649));
nor2 g5823__4547 (.a(n_654), .b(counter_9_), .y(n_644));
nand2 g5824__9682 (.a(n_643), .b(n_178), .y(n_654));
inv g5825 (.a(n_643), .y(n_648));
nor2 g5826__2683 (.a(n_650), .b(counter_7_), .y(n_643));
nand2 g5827__1309 (.a(n_642), .b(n_182), .y(n_650));
inv g5828 (.a(n_642), .y(n_652));
nor2 g5829__6877 (.a(n_655), .b(counter_5_), .y(n_642));
inv g5830 (.a(n_641), .y(n_687));
inv g5831 (.a(n_640), .y(n_717));
inv g5832 (.a(n_639), .y(n_677));
inv g5833 (.a(n_638), .y(n_716));
inv g5834 (.a(n_637), .y(n_715));
inv g5835 (.a(n_636), .y(n_714));
inv g5836 (.a(n_635), .y(n_676));
inv g5837 (.a(n_634), .y(n_713));
inv g5838 (.a(n_633), .y(n_712));
inv g5839 (.a(n_632), .y(n_711));
inv g5840 (.a(n_631), .y(n_675));
inv g5841 (.a(n_630), .y(n_710));
inv g5842 (.a(n_629), .y(n_709));
inv g5843 (.a(n_628), .y(n_708));
inv g5844 (.a(n_627), .y(n_674));
inv g5845 (.a(n_626), .y(n_707));
inv g5846 (.a(n_625), .y(n_718));
inv g5847 (.a(n_624), .y(n_706));
inv g5848 (.a(n_623), .y(n_705));
inv g5849 (.a(n_622), .y(n_673));
inv g5850 (.a(n_621), .y(n_704));
inv g5851 (.a(n_620), .y(n_703));
inv g5852 (.a(n_619), .y(n_702));
inv g5853 (.a(n_618), .y(n_701));
inv g5854 (.a(n_617), .y(n_672));
inv g5855 (.a(n_616), .y(n_700));
inv g5856 (.a(n_615), .y(n_699));
inv g5857 (.a(n_614), .y(n_698));
inv g5858 (.a(n_613), .y(n_686));
inv g5859 (.a(n_612), .y(n_671));
inv g5860 (.a(n_611), .y(n_697));
inv g5861 (.a(n_610), .y(n_696));
nor2 g5862__2900 (.a(n_543), .b(n_527), .y(n_641));
nor2 g5863__2391 (.a(n_572), .b(n_571), .y(n_640));
nor2 g5864__7675 (.a(n_570), .b(n_566), .y(n_639));
nor2 g5865__7118 (.a(n_569), .b(n_568), .y(n_638));
nor2 g5866__8757 (.a(n_567), .b(n_565), .y(n_637));
nor2 g5867__1786 (.a(n_564), .b(n_563), .y(n_636));
nor2 g5868__5953 (.a(n_562), .b(n_558), .y(n_635));
nor2 g5869__5703 (.a(n_561), .b(n_560), .y(n_634));
nor2 g5870__7114 (.a(n_559), .b(n_557), .y(n_633));
nor2 g5871__5266 (.a(n_556), .b(n_555), .y(n_632));
nor2 g5872__2250 (.a(n_554), .b(n_549), .y(n_631));
nor2 g5873__6083 (.a(n_553), .b(n_552), .y(n_630));
nor2 g5874__2703 (.a(n_551), .b(n_550), .y(n_629));
nor2 g5875__5795 (.a(n_548), .b(n_547), .y(n_628));
nor2 g5876__7344 (.a(n_577), .b(n_541), .y(n_627));
nor2 g5877__1840 (.a(n_546), .b(n_544), .y(n_626));
nor2 g5878__5019 (.a(n_574), .b(n_573), .y(n_625));
nor2 g5879__1857 (.a(n_542), .b(n_540), .y(n_624));
nor2 g5880__9906 (.a(n_539), .b(n_538), .y(n_623));
nor2 g5881__8780 (.a(n_536), .b(n_532), .y(n_622));
nor2 g5882__4296 (.a(n_537), .b(n_535), .y(n_621));
nor2 g5883__3772 (.a(n_534), .b(n_533), .y(n_620));
nor2 g5884__1474 (.a(n_531), .b(n_530), .y(n_619));
nor2 g5885__4547 (.a(n_529), .b(n_528), .y(n_618));
nor2 g5886__9682 (.a(n_526), .b(n_523), .y(n_617));
nor2 g5887__2683 (.a(n_525), .b(n_524), .y(n_616));
nor2 g5888__1309 (.a(n_522), .b(n_521), .y(n_615));
nor2 g5889__6877 (.a(n_520), .b(n_519), .y(n_614));
nor2 g5890__2900 (.a(n_515), .b(n_509), .y(n_613));
nor2 g5891__2391 (.a(n_518), .b(n_449), .y(n_612));
nor2 g5892__7675 (.a(n_517), .b(n_516), .y(n_611));
nor2 g5893__7118 (.a(n_514), .b(n_480), .y(n_610));
inv g5894 (.a(n_609), .y(n_683));
inv g5895 (.a(n_608), .y(n_695));
inv g5896 (.a(n_607), .y(n_694));
inv g5897 (.a(n_606), .y(n_693));
inv g5899 (.a(n_604), .y(n_685));
inv g5900 (.a(n_603), .y(n_669));
inv g5904 (.a(n_599), .y(n_668));
inv g5905 (.a(n_598), .y(n_688));
inv g5906 (.a(n_597), .y(n_684));
inv g5907 (.a(n_596), .y(n_667));
inv g5908 (.a(n_595), .y(n_666));
inv g5909 (.a(n_594), .y(n_665));
inv g5910 (.a(n_593), .y(n_670));
inv g5911 (.a(n_592), .y(n_664));
inv g5912 (.a(n_591), .y(n_682));
inv g5913 (.a(n_590), .y(n_663));
inv g5914 (.a(n_589), .y(n_662));
inv g5915 (.a(n_588), .y(n_661));
inv g5916 (.a(n_587), .y(n_681));
inv g5917 (.a(n_586), .y(n_660));
inv g5918 (.a(n_585), .y(n_680));
inv g5919 (.a(n_584), .y(n_659));
inv g5922 (.a(n_581), .y(n_679));
inv g5924 (.a(n_579), .y(n_678));
inv g5925 (.a(n_578), .y(n_719));
nor2 g5926__8757 (.a(n_479), .b(n_476), .y(n_609));
nor2 g5927__1786 (.a(n_511), .b(n_510), .y(n_608));
nor2 g5928__5953 (.a(n_507), .b(n_506), .y(n_607));
nor2 g5929__5703 (.a(n_505), .b(n_504), .y(n_606));
nor2 g5931__5266 (.a(n_497), .b(n_488), .y(n_604));
nor2 g5932__2250 (.a(n_500), .b(n_495), .y(n_603));
nor2 g5936__7344 (.a(n_490), .b(n_487), .y(n_599));
nor2 g5937__1840 (.a(n_491), .b(n_489), .y(n_598));
nor2 g5938__5019 (.a(n_485), .b(n_483), .y(n_597));
nor2 g5939__1857 (.a(n_486), .b(n_484), .y(n_596));
nor2 g5940__9906 (.a(n_482), .b(n_481), .y(n_595));
nor2 g5941__8780 (.a(n_512), .b(n_478), .y(n_594));
nor2 g5942__4296 (.a(n_508), .b(n_503), .y(n_593));
nor2 g5943__3772 (.a(n_477), .b(n_475), .y(n_592));
nor2 g5944__1474 (.a(n_473), .b(n_471), .y(n_591));
nor2 g5945__4547 (.a(n_474), .b(n_472), .y(n_590));
nor2 g5946__9682 (.a(n_470), .b(n_469), .y(n_589));
nor2 g5947__2683 (.a(n_468), .b(n_466), .y(n_588));
nor2 g5948__1309 (.a(n_467), .b(n_464), .y(n_587));
nor2 g5949__6877 (.a(n_465), .b(n_463), .y(n_586));
nor2 g5950__2900 (.a(n_461), .b(n_459), .y(n_585));
nor2 g5951__2391 (.a(n_462), .b(n_460), .y(n_584));
nor2 g5954__8757 (.a(n_455), .b(n_452), .y(n_581));
nor2 g5956__5953 (.a(n_545), .b(n_575), .y(n_579));
nor2 g5957__5703 (.a(n_450), .b(n_576), .y(n_578));
nand2 g5958__7114 (.a(n_3111), .b(n_180), .y(n_655));
nand2 g5959__5266 (.a(n_273), .b(n_308), .y(n_577));
nand2 g5960__2250 (.a(n_349), .b(n_319), .y(n_576));
nand2 g5961__6083 (.a(n_346), .b(n_445), .y(n_575));
nand2 g5962__2703 (.a(n_447), .b(n_347), .y(n_574));
nand2 g5963__5795 (.a(n_345), .b(n_446), .y(n_573));
nand2 g5964__7344 (.a(n_444), .b(n_342), .y(n_572));
nand2 g5965__1840 (.a(n_341), .b(n_443), .y(n_571));
nand2 g5966__5019 (.a(n_339), .b(n_336), .y(n_570));
nand2 g5967__1857 (.a(n_442), .b(n_338), .y(n_569));
nand2 g5968__9906 (.a(n_337), .b(n_441), .y(n_568));
nand2 g5969__8780 (.a(n_440), .b(n_335), .y(n_567));
nand2 g5970__4296 (.a(n_208), .b(n_437), .y(n_566));
nand2 g5971__3772 (.a(n_219), .b(n_439), .y(n_565));
nand2 g5972__1474 (.a(n_436), .b(n_198), .y(n_564));
nand2 g5973__4547 (.a(n_330), .b(n_435), .y(n_563));
nand2 g5974__9682 (.a(n_215), .b(n_325), .y(n_562));
nand2 g5975__2683 (.a(n_434), .b(n_327), .y(n_561));
nand2 g5976__1309 (.a(n_224), .b(n_433), .y(n_560));
nand2 g5977__6877 (.a(n_432), .b(n_324), .y(n_559));
nand2 g5978__2900 (.a(n_230), .b(n_428), .y(n_558));
nand2 g5979__2391 (.a(n_323), .b(n_430), .y(n_557));
nand2 g5980__7675 (.a(n_429), .b(n_321), .y(n_556));
nand2 g5981__7118 (.a(n_241), .b(n_427), .y(n_555));
nand2 g5982__8757 (.a(n_317), .b(n_315), .y(n_554));
nand2 g5983__1786 (.a(n_425), .b(n_318), .y(n_553));
nand2 g5984__5953 (.a(n_316), .b(n_424), .y(n_552));
nand2 g5985__5703 (.a(n_423), .b(n_271), .y(n_551));
nand2 g5986__7114 (.a(n_313), .b(n_422), .y(n_550));
nand2 g5987__5266 (.a(n_312), .b(n_420), .y(n_549));
nand2 g5988__2250 (.a(n_421), .b(n_310), .y(n_548));
nand2 g5989__6083 (.a(n_268), .b(n_419), .y(n_547));
nand2 g5990__2703 (.a(n_418), .b(n_277), .y(n_546));
nand2 g5991__5795 (.a(n_350), .b(n_348), .y(n_545));
nand2 g5992__7344 (.a(n_309), .b(n_416), .y(n_544));
nand2 g5993__1840 (.a(n_307), .b(n_297), .y(n_543));
nand2 g5994__5019 (.a(n_415), .b(n_275), .y(n_542));
nand2 g5995__1857 (.a(n_304), .b(n_409), .y(n_541));
nand2 g5996__9906 (.a(n_306), .b(n_414), .y(n_540));
nand2 g5997__8780 (.a(n_413), .b(n_303), .y(n_539));
nand2 g5998__4296 (.a(n_301), .b(n_411), .y(n_538));
nand2 g5999__3772 (.a(n_410), .b(n_299), .y(n_537));
nand2 g6000__1474 (.a(n_291), .b(n_295), .y(n_536));
nand2 g6001__4547 (.a(n_283), .b(n_408), .y(n_535));
nand2 g6002__9682 (.a(n_407), .b(n_298), .y(n_534));
nand2 g6003__2683 (.a(n_294), .b(n_406), .y(n_533));
nand2 g6004__1309 (.a(n_296), .b(n_404), .y(n_532));
nand2 g6005__6877 (.a(n_405), .b(n_302), .y(n_531));
nand2 g6006__2900 (.a(n_286), .b(n_403), .y(n_530));
nand2 g6007__2391 (.a(n_402), .b(n_288), .y(n_529));
nand2 g6008__7675 (.a(n_193), .b(n_401), .y(n_528));
nand2 g6009__7118 (.a(n_289), .b(n_397), .y(n_527));
nand2 g6010__8757 (.a(n_448), .b(n_331), .y(n_526));
nand2 g6011__1786 (.a(n_399), .b(n_285), .y(n_525));
nand2 g6012__5953 (.a(n_284), .b(n_398), .y(n_524));
nand2 g6013__5703 (.a(n_282), .b(n_394), .y(n_523));
nand2 g6014__7114 (.a(n_431), .b(n_326), .y(n_522));
nand2 g6015__5266 (.a(n_333), .b(n_396), .y(n_521));
nand2 g6016__2250 (.a(n_393), .b(n_328), .y(n_520));
nand2 g6017__6083 (.a(n_352), .b(n_392), .y(n_519));
nand2 g6018__2703 (.a(n_343), .b(n_280), .y(n_518));
nand2 g6019__5795 (.a(n_391), .b(n_340), .y(n_517));
nand2 g6020__7344 (.a(n_249), .b(n_390), .y(n_516));
nand2 g6021__1840 (.a(n_205), .b(n_278), .y(n_515));
nand2 g6022__5019 (.a(n_389), .b(n_196), .y(n_514));
inv g6023 (.a(n_3111), .y(n_646));
nand2 g6024__1857 (.a(n_248), .b(n_247), .y(n_512));
nand2 g6025__9906 (.a(n_387), .b(n_236), .y(n_511));
nand2 g6026__8780 (.a(n_227), .b(n_385), .y(n_510));
nand2 g6027__4296 (.a(n_267), .b(n_412), .y(n_509));
nand2 g6028__3772 (.a(n_255), .b(n_276), .y(n_508));
nand2 g6029__1474 (.a(n_384), .b(n_244), .y(n_507));
nand2 g6030__4547 (.a(n_287), .b(n_383), .y(n_506));
nand2 g6031__9682 (.a(n_382), .b(n_274), .y(n_505));
nand2 g6032__2683 (.a(n_266), .b(n_400), .y(n_504));
nand2 g6033__1309 (.a(n_272), .b(n_426), .y(n_503));
nand2 g6034__6877 (.a(n_381), .b(n_270), .y(n_502));
nand2 g6035__2900 (.a(n_269), .b(n_380), .y(n_501));
nand2 g6036__2391 (.a(n_265), .b(n_320), .y(n_500));
nand2 g6039__8757 (.a(n_264), .b(n_263), .y(n_497));
nand2 g6040__1786 (.a(n_378), .b(n_292), .y(n_496));
nand2 g6041__5953 (.a(n_300), .b(n_376), .y(n_495));
nand2 g6042__5703 (.a(n_305), .b(n_377), .y(n_494));
nand2 g6043__7114 (.a(n_417), .b(n_311), .y(n_493));
nand2 g6044__5266 (.a(n_314), .b(n_438), .y(n_492));
nand2 g6045__2250 (.a(n_375), .b(n_322), .y(n_491));
nand2 g6046__6083 (.a(n_334), .b(n_261), .y(n_490));
nand2 g6047__2703 (.a(n_329), .b(n_374), .y(n_489));
nand2 g6048__5795 (.a(n_260), .b(n_373), .y(n_488));
nand2 g6049__7344 (.a(n_259), .b(n_372), .y(n_487));
nand2 g6050__1840 (.a(n_258), .b(n_257), .y(n_486));
nand2 g6051__5019 (.a(n_256), .b(n_254), .y(n_485));
nand2 g6052__1857 (.a(n_290), .b(n_371), .y(n_484));
nand2 g6053__9906 (.a(n_251), .b(n_369), .y(n_483));
nand2 g6054__8780 (.a(n_253), .b(n_252), .y(n_482));
nand2 g6055__4296 (.a(n_250), .b(n_370), .y(n_481));
nand2 g6056__3772 (.a(n_194), .b(n_388), .y(n_480));
nand2 g6057__1474 (.a(n_246), .b(n_243), .y(n_479));
nand2 g6058__4547 (.a(n_245), .b(n_368), .y(n_478));
nand2 g6059__9682 (.a(n_242), .b(n_240), .y(n_477));
nand2 g6060__2683 (.a(n_239), .b(n_367), .y(n_476));
nand2 g6061__1309 (.a(n_238), .b(n_366), .y(n_475));
nand2 g6062__6877 (.a(n_237), .b(n_235), .y(n_474));
nand2 g6063__2900 (.a(n_234), .b(n_233), .y(n_473));
nand2 g6064__2391 (.a(n_332), .b(n_365), .y(n_472));
nand2 g6065__7675 (.a(n_229), .b(n_363), .y(n_471));
nand2 g6066__7118 (.a(n_232), .b(n_231), .y(n_470));
nand2 g6067__8757 (.a(n_228), .b(n_364), .y(n_469));
nand2 g6068__1786 (.a(n_226), .b(n_225), .y(n_468));
nand2 g6069__5953 (.a(n_223), .b(n_221), .y(n_467));
nand2 g6070__5703 (.a(n_222), .b(n_362), .y(n_466));
nand2 g6071__7114 (.a(n_220), .b(n_218), .y(n_465));
nand2 g6072__5266 (.a(n_217), .b(n_361), .y(n_464));
nand2 g6073__2250 (.a(n_216), .b(n_360), .y(n_463));
nand2 g6074__6083 (.a(n_214), .b(n_213), .y(n_462));
nand2 g6075__2703 (.a(n_212), .b(n_211), .y(n_461));
nand2 g6076__5795 (.a(n_262), .b(n_359), .y(n_460));
nand2 g6077__7344 (.a(n_207), .b(n_357), .y(n_459));
nand2 g6079__5019 (.a(n_206), .b(n_358), .y(n_457));
nand2 g6081__9906 (.a(n_202), .b(n_200), .y(n_455));
nand2 g6084__3772 (.a(n_293), .b(n_355), .y(n_452));
nand2 g6086__4547 (.a(n_353), .b(n_351), .y(n_450));
nand2 g6087__9682 (.a(n_279), .b(n_386), .y(n_449));
nand2 g6089__1309 (.a(n_3841), .b(key_r_80_), .y(n_448));
nand2 g6090__6877 (.a(n_2757), .b(key_r_94_), .y(n_447));
nand2 g6091__2900 (.a(n_191), .b(key_r_126_), .y(n_446));
nand2 g6092__2391 (.a(n_3833), .b(key_r_118_), .y(n_445));
nand2 g6093__7675 (.a(n_2757), .b(key_r_93_), .y(n_444));
nand2 g6094__7118 (.a(n_191), .b(key_r_125_), .y(n_443));
nand2 g6095__8757 (.a(n_2757), .b(key_r_92_), .y(n_442));
nand2 g6096__1786 (.a(n_191), .b(key_r_124_), .y(n_441));
nand2 g6097__5953 (.a(n_2757), .b(key_r_91_), .y(n_440));
nand2 g6098__5703 (.a(n_191), .b(key_r_123_), .y(n_439));
nand2 g6099__7114 (.a(n_191), .b(key_r_97_), .y(n_438));
nand2 g6100__5266 (.a(n_3833), .b(key_r_117_), .y(n_437));
nand2 g6101__2250 (.a(n_2757), .b(key_r_90_), .y(n_436));
nand2 g6102__6083 (.a(n_191), .b(key_r_122_), .y(n_435));
nand2 g6103__2703 (.a(n_2757), .b(key_r_89_), .y(n_434));
nand2 g6104__5795 (.a(n_191), .b(key_r_121_), .y(n_433));
nand2 g6105__7344 (.a(n_2757), .b(key_r_88_), .y(n_432));
nand2 g6106__1840 (.a(n_2757), .b(key_r_75_), .y(n_431));
nand2 g6107__5019 (.a(n_191), .b(key_r_120_), .y(n_430));
nand2 g6108__1857 (.a(n_2757), .b(key_r_87_), .y(n_429));
nand2 g6109__9906 (.a(n_3833), .b(key_r_116_), .y(n_428));
nand2 g6110__8780 (.a(n_191), .b(key_r_119_), .y(n_427));
nand2 g6111__4296 (.a(n_3833), .b(key_r_110_), .y(n_426));
nand2 g6112__3772 (.a(n_2757), .b(key_r_86_), .y(n_425));
nand2 g6113__1474 (.a(n_191), .b(key_r_118_), .y(n_424));
nand2 g6114__4547 (.a(n_2757), .b(key_r_85_), .y(n_423));
nand2 g6115__9682 (.a(n_191), .b(key_r_117_), .y(n_422));
nand2 g6116__2683 (.a(n_2757), .b(key_r_84_), .y(n_421));
nand2 g6117__1309 (.a(n_3833), .b(key_r_115_), .y(n_420));
nand2 g6118__6877 (.a(n_191), .b(key_r_116_), .y(n_419));
nand2 g6119__2900 (.a(n_2757), .b(key_r_83_), .y(n_418));
nand2 g6120__2391 (.a(n_2757), .b(key_r_65_), .y(n_417));
nand2 g6121__7675 (.a(n_191), .b(key_r_115_), .y(n_416));
nand2 g6122__7118 (.a(n_2757), .b(key_r_82_), .y(n_415));
nand2 g6123__8757 (.a(n_191), .b(key_r_114_), .y(n_414));
nand2 g6124__1786 (.a(n_2757), .b(key_r_81_), .y(n_413));
nand2 g6125__5953 (.a(n_3833), .b(key_r_126_), .y(n_412));
nand2 g6126__5703 (.a(n_191), .b(key_r_113_), .y(n_411));
nand2 g6127__7114 (.a(n_2757), .b(key_r_80_), .y(n_410));
nand2 g6128__5266 (.a(n_3833), .b(key_r_114_), .y(n_409));
nand2 g6129__2250 (.a(n_191), .b(key_r_112_), .y(n_408));
nand2 g6130__6083 (.a(n_2757), .b(key_r_79_), .y(n_407));
nand2 g6131__2703 (.a(n_191), .b(key_r_111_), .y(n_406));
nand2 g6132__5795 (.a(n_2757), .b(key_r_78_), .y(n_405));
nand2 g6133__7344 (.a(n_3833), .b(key_r_113_), .y(n_404));
nand2 g6134__1840 (.a(n_191), .b(key_r_110_), .y(n_403));
nand2 g6135__5019 (.a(n_2757), .b(key_r_77_), .y(n_402));
nand2 g6136__1857 (.a(n_191), .b(key_r_109_), .y(n_401));
nand2 g6137__9906 (.a(n_191), .b(key_r_101_), .y(n_400));
nand2 g6138__8780 (.a(n_2757), .b(key_r_76_), .y(n_399));
nand2 g6139__4296 (.a(n_191), .b(key_r_108_), .y(n_398));
nand2 g6140__3772 (.a(n_3833), .b(key_r_127_), .y(n_397));
nand2 g6141__1474 (.a(n_191), .b(key_r_107_), .y(n_396));
nand2 g6142__4547 (.a(n_2757), .b(key_r_67_), .y(n_395));
nand2 g6143__9682 (.a(n_3833), .b(key_r_112_), .y(n_394));
nand2 g6144__2683 (.a(n_2757), .b(key_r_74_), .y(n_393));
nand2 g6145__1309 (.a(n_191), .b(key_r_106_), .y(n_392));
nand2 g6146__6877 (.a(n_2757), .b(key_r_73_), .y(n_391));
nand2 g6147__2900 (.a(n_191), .b(key_r_105_), .y(n_390));
nand2 g6148__2391 (.a(n_2757), .b(key_r_72_), .y(n_389));
nand2 g6149__7675 (.a(n_191), .b(key_r_104_), .y(n_388));
nand2 g6150__7118 (.a(n_2757), .b(key_r_71_), .y(n_387));
nand2 g6151__8757 (.a(n_3833), .b(key_r_111_), .y(n_386));
nand2 g6152__1786 (.a(n_191), .b(key_r_103_), .y(n_385));
nand2 g6153__5953 (.a(n_2757), .b(key_r_70_), .y(n_384));
nand2 g6154__5703 (.a(n_191), .b(key_r_102_), .y(n_383));
nand2 g6155__7114 (.a(n_2757), .b(key_r_69_), .y(n_382));
nand2 g6156__5266 (.a(n_2757), .b(key_r_68_), .y(n_381));
nand2 g6157__2250 (.a(n_191), .b(key_r_100_), .y(n_380));
nand2 g6158__6083 (.a(n_191), .b(key_r_99_), .y(n_379));
nand2 g6159__2703 (.a(n_2757), .b(key_r_66_), .y(n_378));
nand2 g6160__5795 (.a(n_191), .b(key_r_98_), .y(n_377));
nand2 g6161__7344 (.a(n_3833), .b(key_r_109_), .y(n_376));
nand2 g6162__1840 (.a(n_2757), .b(key_r_64_), .y(n_375));
nand2 g6163__5019 (.a(n_191), .b(key_r_96_), .y(n_374));
nand2 g6164__1857 (.a(n_3833), .b(key_r_125_), .y(n_373));
nand2 g6165__9906 (.a(n_3833), .b(key_r_108_), .y(n_372));
nand2 g6166__8780 (.a(n_3833), .b(key_r_107_), .y(n_371));
nand2 g6167__4296 (.a(n_3833), .b(key_r_106_), .y(n_370));
nand2 g6168__3772 (.a(n_3833), .b(key_r_124_), .y(n_369));
nand2 g6169__1474 (.a(n_3833), .b(key_r_105_), .y(n_368));
nand2 g6170__4547 (.a(n_3833), .b(key_r_123_), .y(n_367));
nand2 g6171__9682 (.a(n_3833), .b(key_r_104_), .y(n_366));
nand2 g6172__2683 (.a(n_3833), .b(key_r_103_), .y(n_365));
nand2 g6173__1309 (.a(n_3833), .b(key_r_102_), .y(n_364));
nand2 g6174__6877 (.a(n_3833), .b(key_r_122_), .y(n_363));
nand2 g6175__2900 (.a(n_3833), .b(key_r_101_), .y(n_362));
nand2 g6176__2391 (.a(n_3833), .b(key_r_121_), .y(n_361));
nand2 g6177__7675 (.a(n_3833), .b(key_r_100_), .y(n_360));
nand2 g6178__7118 (.a(n_3833), .b(key_r_99_), .y(n_359));
nand2 g6179__8757 (.a(n_3833), .b(key_r_98_), .y(n_358));
nand2 g6180__1786 (.a(n_3833), .b(key_r_120_), .y(n_357));
nand2 g6182__5703 (.a(n_3833), .b(key_r_119_), .y(n_355));
nand2 g6184__5266 (.a(n_2757), .b(key_r_95_), .y(n_353));
nand2 g6185__2250 (.a(n_2758), .b(key_r_10_), .y(n_352));
nand2 g6186__6083 (.a(n_187), .b(key_r_63_), .y(n_351));
nand2 g6187__2703 (.a(n_3841), .b(key_r_86_), .y(n_350));
nand2 g6188__5795 (.a(n_2758), .b(key_r_31_), .y(n_349));
nand2 g6189__7344 (.a(n_3842), .b(key_r_54_), .y(n_348));
nand2 g6190__1840 (.a(n_187), .b(key_r_62_), .y(n_347));
nand2 g6191__5019 (.a(n_3832), .b(key_r_22_), .y(n_346));
nand2 g6192__1857 (.a(n_2758), .b(key_r_30_), .y(n_345));
nand2 g6193__9906 (.a(n_2758), .b(key_r_3_), .y(n_344));
nand2 g6194__8780 (.a(n_3841), .b(key_r_79_), .y(n_343));
nand2 g6195__4296 (.a(n_187), .b(key_r_61_), .y(n_342));
nand2 g6196__3772 (.a(n_2758), .b(key_r_29_), .y(n_341));
nand2 g6197__1474 (.a(n_187), .b(key_r_41_), .y(n_340));
nand2 g6198__4547 (.a(n_3841), .b(key_r_85_), .y(n_339));
nand2 g6199__9682 (.a(n_187), .b(key_r_60_), .y(n_338));
nand2 g6200__2683 (.a(n_2758), .b(key_r_28_), .y(n_337));
nand2 g6201__1309 (.a(n_3842), .b(key_r_53_), .y(n_336));
nand2 g6202__6877 (.a(n_187), .b(key_r_59_), .y(n_335));
nand2 g6203__2900 (.a(n_3841), .b(key_r_76_), .y(n_334));
nand2 g6204__2391 (.a(n_2758), .b(key_r_11_), .y(n_333));
nand2 g6205__7675 (.a(n_3832), .b(key_r_7_), .y(n_332));
nand2 g6206__7118 (.a(n_3842), .b(key_r_48_), .y(n_331));
nand2 g6207__8757 (.a(n_2758), .b(key_r_26_), .y(n_330));
nand2 g6208__1786 (.a(n_2758), .b(key_r_0_), .y(n_329));
nand2 g6209__5953 (.a(n_187), .b(key_r_42_), .y(n_328));
nand2 g6210__5703 (.a(n_187), .b(key_r_57_), .y(n_327));
nand2 g6211__7114 (.a(n_187), .b(key_r_43_), .y(n_326));
nand2 g6212__5266 (.a(n_3842), .b(key_r_52_), .y(n_325));
nand2 g6213__2250 (.a(n_187), .b(key_r_56_), .y(n_324));
nand2 g6214__6083 (.a(n_2758), .b(key_r_24_), .y(n_323));
nand2 g6215__2703 (.a(n_187), .b(key_r_32_), .y(n_322));
nand2 g6216__5795 (.a(n_187), .b(key_r_55_), .y(n_321));
nand2 g6217__7344 (.a(n_3842), .b(key_r_45_), .y(n_320));
nand2 g6218__1840 (.a(n_191), .b(key_r_127_), .y(n_319));
nand2 g6219__5019 (.a(n_187), .b(key_r_54_), .y(n_318));
nand2 g6220__1857 (.a(n_3841), .b(key_r_83_), .y(n_317));
nand2 g6221__9906 (.a(n_2758), .b(key_r_22_), .y(n_316));
nand2 g6222__8780 (.a(n_3842), .b(key_r_51_), .y(n_315));
nand2 g6223__4296 (.a(n_2758), .b(key_r_1_), .y(n_314));
nand2 g6224__3772 (.a(n_2758), .b(key_r_21_), .y(n_313));
nand2 g6225__1474 (.a(n_3832), .b(key_r_19_), .y(n_312));
nand2 g6226__4547 (.a(n_187), .b(key_r_33_), .y(n_311));
nand2 g6227__9682 (.a(n_187), .b(key_r_52_), .y(n_310));
xor2 g6229__1309 (.a(v1_22_), .b(v1_13_), .y(n_953));
nand2 g6230__6877 (.a(n_2758), .b(key_r_19_), .y(n_309));
nand2 g6231__2900 (.a(n_3842), .b(key_r_50_), .y(n_308));
nand2 g6232__2391 (.a(n_3841), .b(key_r_95_), .y(n_307));
nand2 g6233__7675 (.a(n_2758), .b(key_r_18_), .y(n_306));
nand2 g6234__7118 (.a(n_2758), .b(key_r_2_), .y(n_305));
nand2 g6235__8757 (.a(n_3832), .b(key_r_18_), .y(n_304));
nand2 g6236__1786 (.a(n_187), .b(key_r_49_), .y(n_303));
nand2 g6237__5953 (.a(n_187), .b(key_r_46_), .y(n_302));
nand2 g6238__5703 (.a(n_2758), .b(key_r_17_), .y(n_301));
nand2 g6239__7114 (.a(n_3832), .b(key_r_13_), .y(n_300));
nand2 g6240__5266 (.a(n_187), .b(key_r_48_), .y(n_299));
nand2 g6241__2250 (.a(n_187), .b(key_r_47_), .y(n_298));
nand2 g6242__6083 (.a(n_3842), .b(key_r_63_), .y(n_297));
nand2 g6243__2703 (.a(n_3832), .b(key_r_17_), .y(n_296));
nand2 g6244__5795 (.a(n_3842), .b(key_r_49_), .y(n_295));
nand2 g6245__7344 (.a(n_2758), .b(key_r_15_), .y(n_294));
nand2 g6246__1840 (.a(n_3832), .b(key_r_23_), .y(n_293));
nand2 g6247__5019 (.a(n_187), .b(key_r_34_), .y(n_292));
nand2 g6248__1857 (.a(n_3841), .b(key_r_81_), .y(n_291));
nand2 g6249__9906 (.a(n_3832), .b(key_r_11_), .y(n_290));
nand2 g6250__8780 (.a(n_3832), .b(key_r_31_), .y(n_289));
nand2 g6251__4296 (.a(n_187), .b(key_r_45_), .y(n_288));
nand2 g6252__3772 (.a(n_2758), .b(key_r_6_), .y(n_287));
nand2 g6253__1474 (.a(n_2758), .b(key_r_14_), .y(n_286));
nand2 g6254__4547 (.a(n_187), .b(key_r_44_), .y(n_285));
nand2 g6255__9682 (.a(n_2758), .b(key_r_12_), .y(n_284));
nand2 g6256__2683 (.a(n_2758), .b(key_r_16_), .y(n_283));
nand2 g6257__1309 (.a(n_3832), .b(key_r_16_), .y(n_282));
nand2 g6258__6877 (.a(n_187), .b(key_r_35_), .y(n_281));
nand2 g6259__2900 (.a(n_3842), .b(key_r_47_), .y(n_280));
nand2 g6260__2391 (.a(n_3832), .b(key_r_15_), .y(n_279));
nand2 g6261__7675 (.a(n_3842), .b(key_r_62_), .y(n_278));
nand2 g6262__7118 (.a(n_187), .b(key_r_51_), .y(n_277));
nand2 g6263__8757 (.a(n_3842), .b(key_r_46_), .y(n_276));
nand2 g6264__1786 (.a(n_187), .b(key_r_50_), .y(n_275));
nand2 g6265__5953 (.a(n_187), .b(key_r_37_), .y(n_274));
nand2 g6266__5703 (.a(n_3841), .b(key_r_82_), .y(n_273));
nand2 g6267__7114 (.a(n_3832), .b(key_r_14_), .y(n_272));
nand2 g6268__5266 (.a(n_187), .b(key_r_53_), .y(n_271));
nand2 g6269__2250 (.a(n_187), .b(key_r_36_), .y(n_270));
nand2 g6270__6083 (.a(n_2758), .b(key_r_4_), .y(n_269));
nand2 g6271__2703 (.a(n_2758), .b(key_r_20_), .y(n_268));
nand2 g6272__5795 (.a(n_3832), .b(key_r_30_), .y(n_267));
nand2 g6273__7344 (.a(n_2758), .b(key_r_5_), .y(n_266));
nand2 g6274__1840 (.a(n_3841), .b(key_r_77_), .y(n_265));
nand2 g6275__5019 (.a(n_3841), .b(key_r_93_), .y(n_264));
nand2 g6276__1857 (.a(n_3842), .b(key_r_61_), .y(n_263));
nand2 g6277__9906 (.a(n_3832), .b(key_r_3_), .y(n_262));
nand2 g6278__8780 (.a(n_3842), .b(key_r_44_), .y(n_261));
nand2 g6279__4296 (.a(n_3832), .b(key_r_29_), .y(n_260));
nand2 g6280__3772 (.a(n_3832), .b(key_r_12_), .y(n_259));
nand2 g6281__1474 (.a(n_3841), .b(key_r_75_), .y(n_258));
nand2 g6282__4547 (.a(n_3842), .b(key_r_43_), .y(n_257));
nand2 g6283__9682 (.a(n_3841), .b(key_r_92_), .y(n_256));
nand2 g6284__2683 (.a(n_3841), .b(key_r_78_), .y(n_255));
nand2 g6285__1309 (.a(n_3842), .b(key_r_60_), .y(n_254));
nand2 g6286__6877 (.a(n_3841), .b(key_r_74_), .y(n_253));
nand2 g6287__2900 (.a(n_3842), .b(key_r_42_), .y(n_252));
nand2 g6288__2391 (.a(n_3832), .b(key_r_28_), .y(n_251));
nand2 g6289__7675 (.a(n_3832), .b(key_r_10_), .y(n_250));
nand2 g6290__7118 (.a(n_2758), .b(key_r_9_), .y(n_249));
nand2 g6291__8757 (.a(n_3841), .b(key_r_73_), .y(n_248));
nand2 g6292__1786 (.a(n_3842), .b(key_r_41_), .y(n_247));
nand2 g6293__5953 (.a(n_3841), .b(key_r_91_), .y(n_246));
nand2 g6294__5703 (.a(n_3832), .b(key_r_9_), .y(n_245));
nand2 g6295__7114 (.a(n_187), .b(key_r_38_), .y(n_244));
nand2 g6296__5266 (.a(n_3842), .b(key_r_59_), .y(n_243));
nand2 g6297__2250 (.a(n_3841), .b(key_r_72_), .y(n_242));
nand2 g6298__6083 (.a(n_2758), .b(key_r_23_), .y(n_241));
nand2 g6299__2703 (.a(n_3842), .b(key_r_40_), .y(n_240));
nand2 g6300__5795 (.a(n_3832), .b(key_r_27_), .y(n_239));
nand2 g6301__7344 (.a(n_3832), .b(key_r_8_), .y(n_238));
nand2 g6302__1840 (.a(n_3841), .b(key_r_71_), .y(n_237));
nand2 g6303__5019 (.a(n_187), .b(key_r_39_), .y(n_236));
nand2 g6304__1857 (.a(n_3842), .b(key_r_39_), .y(n_235));
nand2 g6305__9906 (.a(n_3841), .b(key_r_90_), .y(n_234));
nand2 g6306__8780 (.a(n_3842), .b(key_r_58_), .y(n_233));
nand2 g6307__4296 (.a(n_3841), .b(key_r_70_), .y(n_232));
nand2 g6308__3772 (.a(n_3842), .b(key_r_38_), .y(n_231));
nand2 g6309__1474 (.a(n_3832), .b(key_r_20_), .y(n_230));
nand2 g6310__4547 (.a(n_3832), .b(key_r_26_), .y(n_229));
nand2 g6311__9682 (.a(n_3832), .b(key_r_6_), .y(n_228));
nand2 g6312__2683 (.a(n_2758), .b(key_r_7_), .y(n_227));
nand2 g6313__1309 (.a(n_3841), .b(key_r_69_), .y(n_226));
nand2 g6314__6877 (.a(n_3842), .b(key_r_37_), .y(n_225));
nand2 g6315__2900 (.a(n_2758), .b(key_r_25_), .y(n_224));
nand2 g6316__2391 (.a(n_3841), .b(key_r_89_), .y(n_223));
nand2 g6317__7675 (.a(n_3832), .b(key_r_5_), .y(n_222));
nand2 g6318__7118 (.a(n_3842), .b(key_r_57_), .y(n_221));
nand2 g6319__8757 (.a(n_3841), .b(key_r_68_), .y(n_220));
nand2 g6320__1786 (.a(n_2758), .b(key_r_27_), .y(n_219));
nand2 g6321__5953 (.a(n_3842), .b(key_r_36_), .y(n_218));
nand2 g6322__5703 (.a(n_3832), .b(key_r_25_), .y(n_217));
nand2 g6323__7114 (.a(n_3832), .b(key_r_4_), .y(n_216));
nand2 g6324__5266 (.a(n_3841), .b(key_r_84_), .y(n_215));
nand2 g6325__2250 (.a(n_3841), .b(key_r_67_), .y(n_214));
nand2 g6326__6083 (.a(n_3842), .b(key_r_35_), .y(n_213));
nand2 g6327__2703 (.a(n_3841), .b(key_r_88_), .y(n_212));
nand2 g6328__5795 (.a(n_3842), .b(key_r_56_), .y(n_211));
nand2 g6331__5019 (.a(n_3832), .b(key_r_21_), .y(n_208));
nand2 g6332__1857 (.a(n_3832), .b(key_r_24_), .y(n_207));
nand2 g6333__9906 (.a(n_3832), .b(key_r_2_), .y(n_206));
nand2 g6334__8780 (.a(n_3841), .b(key_r_94_), .y(n_205));
nand2 g6337__1474 (.a(n_3841), .b(key_r_87_), .y(n_202));
nand2 g6339__9682 (.a(n_3842), .b(key_r_55_), .y(n_200));
nand2 g6341__1309 (.a(n_187), .b(key_r_58_), .y(n_198));
nand2 g6343__2900 (.a(n_187), .b(key_r_40_), .y(n_196));
nand2 g6345__7675 (.a(n_2758), .b(key_r_8_), .y(n_194));
xor2 g6346__7118 (.a(v1_31_), .b(v1_22_), .y(n_944));
xor2 g6347__8757 (.a(v1_17_), .b(v1_8_), .y(n_958));
xor2 g6348__1786 (.a(v1_9_), .b(v1_0_), .y(n_966));
xor2 g6349__5953 (.a(v1_13_), .b(v1_4_), .y(n_962));
xor2 g6350__5703 (.a(v1_29_), .b(v1_20_), .y(n_946));
xor2 g6351__7114 (.a(v1_30_), .b(v1_21_), .y(n_945));
xor2 g6352__5266 (.a(v1_28_), .b(v1_19_), .y(n_947));
xor2 g6353__2250 (.a(v1_27_), .b(v1_18_), .y(n_948));
xor2 g6354__6083 (.a(v1_26_), .b(v1_17_), .y(n_949));
xor2 g6355__2703 (.a(v1_25_), .b(v1_16_), .y(n_950));
xor2 g6356__5795 (.a(v1_24_), .b(v1_15_), .y(n_951));
xor2 g6357__7344 (.a(v1_23_), .b(v1_14_), .y(n_952));
xor2 g6358__1840 (.a(v1_20_), .b(v1_11_), .y(n_955));
xor2 g6359__5019 (.a(v1_19_), .b(v1_10_), .y(n_956));
xor2 g6360__1857 (.a(v1_18_), .b(v1_9_), .y(n_957));
xor2 g6361__9906 (.a(v1_16_), .b(v1_7_), .y(n_959));
xor2 g6362__8780 (.a(v1_15_), .b(v1_6_), .y(n_960));
xor2 g6363__4296 (.a(v1_14_), .b(v1_5_), .y(n_961));
xor2 g6364__3772 (.a(v1_12_), .b(v1_3_), .y(n_963));
xor2 g6365__1474 (.a(v1_11_), .b(v1_2_), .y(n_964));
xor2 g6366__4547 (.a(v1_21_), .b(v1_12_), .y(n_954));
xor2 g6367__9682 (.a(v1_10_), .b(v1_1_), .y(n_965));
nand2 g6368__2683 (.a(n_2758), .b(key_r_13_), .y(n_193));
inv g6369 (.a(n_192), .y(n_653));
nor2 g6370__1309 (.a(counter_1_), .b(sum_0_), .y(n_192));
nor2 g6371__6877 (.a(sum_1_), .b(sum_0_), .y(n_191));
nor2 g6376__7118 (.a(n_179), .b(sum_0_), .y(n_187));
inv g6380 (.a(counter_6_), .y(n_182));
inv g6381 (.a(counter_2_), .y(n_181));
inv g6382 (.a(counter_4_), .y(n_180));
inv g6383 (.a(sum_1_), .y(n_179));
inv g6384 (.a(counter_8_), .y(n_178));
dffr counter_reg_0_ (.rb(reset), .ck(clk), .d(n_80), .q(sum_0_));
dffr counter_reg_1_ (.rb(reset), .ck(clk), .d(n_173), .q(counter_1_));
dffr counter_reg_2_ (.rb(reset), .ck(clk), .d(n_172), .q(counter_2_));
dffr counter_reg_3_ (.rb(reset), .ck(clk), .d(n_170), .q(counter_3_));
dffr counter_reg_4_ (.rb(reset), .ck(clk), .d(n_171), .q(counter_4_));
dffs counter_reg_5_ (.sb(reset), .ck(clk), .d(n_0), .q(counter_5_));
dffr counter_reg_6_ (.rb(reset), .ck(clk), .d(n_168), .q(counter_6_));
dffr counter_reg_7_ (.rb(reset), .ck(clk), .d(n_169), .q(counter_7_));
dffr counter_reg_8_ (.rb(reset), .ck(clk), .d(n_167), .q(counter_8_));
dffr counter_reg_9_ (.rb(reset), .ck(clk), .d(n_166), .q(counter_9_));
dffr counter_reg_10_ (.rb(reset), .ck(clk), .d(n_165), .q(counter_10_));
dffenr key_r_reg_0_ (.rb(reset), .ck(clk), .d(key_0), .en(n_48), .q(key_r_0_));
dffenr key_r_reg_1_ (.rb(reset), .ck(clk), .d(key_1), .en(n_48), .q(key_r_1_));
dffenr key_r_reg_2_ (.rb(reset), .ck(clk), .d(key_2), .en(n_48), .q(key_r_2_));
dffenr key_r_reg_3_ (.rb(reset), .ck(clk), .d(key_3), .en(n_48), .q(key_r_3_));
dffenr key_r_reg_4_ (.rb(reset), .ck(clk), .d(key_4), .en(n_48), .q(key_r_4_));
dffenr key_r_reg_5_ (.rb(reset), .ck(clk), .d(key_5), .en(n_48), .q(key_r_5_));
dffenr key_r_reg_6_ (.rb(reset), .ck(clk), .d(key_6), .en(n_48), .q(key_r_6_));
dffenr key_r_reg_7_ (.rb(reset), .ck(clk), .d(key_7), .en(n_48), .q(key_r_7_));
dffenr key_r_reg_8_ (.rb(reset), .ck(clk), .d(key_8), .en(n_48), .q(key_r_8_));
dffenr key_r_reg_9_ (.rb(reset), .ck(clk), .d(key_9), .en(n_48), .q(key_r_9_));
dffenr key_r_reg_10_ (.rb(reset), .ck(clk), .d(key_10), .en(n_48), .q(key_r_10_));
dffenr key_r_reg_11_ (.rb(reset), .ck(clk), .d(key_11), .en(n_48), .q(key_r_11_));
dffenr key_r_reg_12_ (.rb(reset), .ck(clk), .d(key_12), .en(n_48), .q(key_r_12_));
dffenr key_r_reg_13_ (.rb(reset), .ck(clk), .d(key_13), .en(n_48), .q(key_r_13_));
dffenr key_r_reg_14_ (.rb(reset), .ck(clk), .d(key_14), .en(n_48), .q(key_r_14_));
dffenr key_r_reg_15_ (.rb(reset), .ck(clk), .d(key_15), .en(n_48), .q(key_r_15_));
dffenr key_r_reg_16_ (.rb(reset), .ck(clk), .d(key_16), .en(n_48), .q(key_r_16_));
dffenr key_r_reg_17_ (.rb(reset), .ck(clk), .d(key_17), .en(n_48), .q(key_r_17_));
dffenr key_r_reg_18_ (.rb(reset), .ck(clk), .d(key_18), .en(n_48), .q(key_r_18_));
dffenr key_r_reg_19_ (.rb(reset), .ck(clk), .d(key_19), .en(n_48), .q(key_r_19_));
dffenr key_r_reg_20_ (.rb(reset), .ck(clk), .d(key_20), .en(n_48), .q(key_r_20_));
dffenr key_r_reg_21_ (.rb(reset), .ck(clk), .d(key_21), .en(n_48), .q(key_r_21_));
dffenr key_r_reg_22_ (.rb(reset), .ck(clk), .d(key_22), .en(n_48), .q(key_r_22_));
dffenr key_r_reg_23_ (.rb(reset), .ck(clk), .d(key_23), .en(n_48), .q(key_r_23_));
dffenr key_r_reg_24_ (.rb(reset), .ck(clk), .d(key_24), .en(n_48), .q(key_r_24_));
dffenr key_r_reg_25_ (.rb(reset), .ck(clk), .d(key_25), .en(n_48), .q(key_r_25_));
dffenr key_r_reg_26_ (.rb(reset), .ck(clk), .d(key_26), .en(n_48), .q(key_r_26_));
dffenr key_r_reg_27_ (.rb(reset), .ck(clk), .d(key_27), .en(n_48), .q(key_r_27_));
dffenr key_r_reg_28_ (.rb(reset), .ck(clk), .d(key_28), .en(n_48), .q(key_r_28_));
dffenr key_r_reg_29_ (.rb(reset), .ck(clk), .d(key_29), .en(n_48), .q(key_r_29_));
dffenr key_r_reg_30_ (.rb(reset), .ck(clk), .d(key_30), .en(n_48), .q(key_r_30_));
dffenr key_r_reg_31_ (.rb(reset), .ck(clk), .d(key_31), .en(n_48), .q(key_r_31_));
dffenr key_r_reg_32_ (.rb(reset), .ck(clk), .d(key_32), .en(n_48), .q(key_r_32_));
dffenr key_r_reg_33_ (.rb(reset), .ck(clk), .d(key_33), .en(n_48), .q(key_r_33_));
dffenr key_r_reg_34_ (.rb(reset), .ck(clk), .d(key_34), .en(n_48), .q(key_r_34_));
dffenr key_r_reg_35_ (.rb(reset), .ck(clk), .d(key_35), .en(n_48), .q(key_r_35_));
dffenr key_r_reg_36_ (.rb(reset), .ck(clk), .d(key_36), .en(n_48), .q(key_r_36_));
dffenr key_r_reg_37_ (.rb(reset), .ck(clk), .d(key_37), .en(n_48), .q(key_r_37_));
dffenr key_r_reg_38_ (.rb(reset), .ck(clk), .d(key_38), .en(n_48), .q(key_r_38_));
dffenr key_r_reg_39_ (.rb(reset), .ck(clk), .d(key_39), .en(n_48), .q(key_r_39_));
dffenr key_r_reg_40_ (.rb(reset), .ck(clk), .d(key_40), .en(n_48), .q(key_r_40_));
dffenr key_r_reg_41_ (.rb(reset), .ck(clk), .d(key_41), .en(n_48), .q(key_r_41_));
dffenr key_r_reg_42_ (.rb(reset), .ck(clk), .d(key_42), .en(n_48), .q(key_r_42_));
dffenr key_r_reg_43_ (.rb(reset), .ck(clk), .d(key_43), .en(n_48), .q(key_r_43_));
dffenr key_r_reg_44_ (.rb(reset), .ck(clk), .d(key_44), .en(n_48), .q(key_r_44_));
dffenr key_r_reg_45_ (.rb(reset), .ck(clk), .d(key_45), .en(n_48), .q(key_r_45_));
dffenr key_r_reg_46_ (.rb(reset), .ck(clk), .d(key_46), .en(n_48), .q(key_r_46_));
dffenr key_r_reg_47_ (.rb(reset), .ck(clk), .d(key_47), .en(n_48), .q(key_r_47_));
dffenr key_r_reg_48_ (.rb(reset), .ck(clk), .d(key_48), .en(n_48), .q(key_r_48_));
dffenr key_r_reg_49_ (.rb(reset), .ck(clk), .d(key_49), .en(n_48), .q(key_r_49_));
dffenr key_r_reg_50_ (.rb(reset), .ck(clk), .d(key_50), .en(n_48), .q(key_r_50_));
dffenr key_r_reg_51_ (.rb(reset), .ck(clk), .d(key_51), .en(n_48), .q(key_r_51_));
dffenr key_r_reg_52_ (.rb(reset), .ck(clk), .d(key_52), .en(n_48), .q(key_r_52_));
dffenr key_r_reg_53_ (.rb(reset), .ck(clk), .d(key_53), .en(n_48), .q(key_r_53_));
dffenr key_r_reg_54_ (.rb(reset), .ck(clk), .d(key_54), .en(n_48), .q(key_r_54_));
dffenr key_r_reg_55_ (.rb(reset), .ck(clk), .d(key_55), .en(n_48), .q(key_r_55_));
dffenr key_r_reg_56_ (.rb(reset), .ck(clk), .d(key_56), .en(n_48), .q(key_r_56_));
dffenr key_r_reg_57_ (.rb(reset), .ck(clk), .d(key_57), .en(n_48), .q(key_r_57_));
dffenr key_r_reg_58_ (.rb(reset), .ck(clk), .d(key_58), .en(n_48), .q(key_r_58_));
dffenr key_r_reg_59_ (.rb(reset), .ck(clk), .d(key_59), .en(n_48), .q(key_r_59_));
dffenr key_r_reg_60_ (.rb(reset), .ck(clk), .d(key_60), .en(n_48), .q(key_r_60_));
dffenr key_r_reg_61_ (.rb(reset), .ck(clk), .d(key_61), .en(n_48), .q(key_r_61_));
dffenr key_r_reg_62_ (.rb(reset), .ck(clk), .d(key_62), .en(n_48), .q(key_r_62_));
dffenr key_r_reg_63_ (.rb(reset), .ck(clk), .d(key_63), .en(n_48), .q(key_r_63_));
dffenr key_r_reg_64_ (.rb(reset), .ck(clk), .d(key_64), .en(n_48), .q(key_r_64_));
dffenr key_r_reg_65_ (.rb(reset), .ck(clk), .d(key_65), .en(n_48), .q(key_r_65_));
dffenr key_r_reg_66_ (.rb(reset), .ck(clk), .d(key_66), .en(n_48), .q(key_r_66_));
dffenr key_r_reg_67_ (.rb(reset), .ck(clk), .d(key_67), .en(n_48), .q(key_r_67_));
dffenr key_r_reg_68_ (.rb(reset), .ck(clk), .d(key_68), .en(n_48), .q(key_r_68_));
dffenr key_r_reg_69_ (.rb(reset), .ck(clk), .d(key_69), .en(n_48), .q(key_r_69_));
dffenr key_r_reg_70_ (.rb(reset), .ck(clk), .d(key_70), .en(n_48), .q(key_r_70_));
dffenr key_r_reg_71_ (.rb(reset), .ck(clk), .d(key_71), .en(n_48), .q(key_r_71_));
dffenr key_r_reg_72_ (.rb(reset), .ck(clk), .d(key_72), .en(n_48), .q(key_r_72_));
dffenr key_r_reg_73_ (.rb(reset), .ck(clk), .d(key_73), .en(n_48), .q(key_r_73_));
dffenr key_r_reg_74_ (.rb(reset), .ck(clk), .d(key_74), .en(n_48), .q(key_r_74_));
dffenr key_r_reg_75_ (.rb(reset), .ck(clk), .d(key_75), .en(n_48), .q(key_r_75_));
dffenr key_r_reg_76_ (.rb(reset), .ck(clk), .d(key_76), .en(n_48), .q(key_r_76_));
dffenr key_r_reg_77_ (.rb(reset), .ck(clk), .d(key_77), .en(n_48), .q(key_r_77_));
dffenr key_r_reg_78_ (.rb(reset), .ck(clk), .d(key_78), .en(n_48), .q(key_r_78_));
dffenr key_r_reg_79_ (.rb(reset), .ck(clk), .d(key_79), .en(n_48), .q(key_r_79_));
dffenr key_r_reg_80_ (.rb(reset), .ck(clk), .d(key_80), .en(n_48), .q(key_r_80_));
dffenr key_r_reg_81_ (.rb(reset), .ck(clk), .d(key_81), .en(n_48), .q(key_r_81_));
dffenr key_r_reg_82_ (.rb(reset), .ck(clk), .d(key_82), .en(n_48), .q(key_r_82_));
dffenr key_r_reg_83_ (.rb(reset), .ck(clk), .d(key_83), .en(n_48), .q(key_r_83_));
dffenr key_r_reg_84_ (.rb(reset), .ck(clk), .d(key_84), .en(n_48), .q(key_r_84_));
dffenr key_r_reg_85_ (.rb(reset), .ck(clk), .d(key_85), .en(n_48), .q(key_r_85_));
dffenr key_r_reg_86_ (.rb(reset), .ck(clk), .d(key_86), .en(n_48), .q(key_r_86_));
dffenr key_r_reg_87_ (.rb(reset), .ck(clk), .d(key_87), .en(n_48), .q(key_r_87_));
dffenr key_r_reg_88_ (.rb(reset), .ck(clk), .d(key_88), .en(n_48), .q(key_r_88_));
dffenr key_r_reg_89_ (.rb(reset), .ck(clk), .d(key_89), .en(n_48), .q(key_r_89_));
dffenr key_r_reg_90_ (.rb(reset), .ck(clk), .d(key_90), .en(n_48), .q(key_r_90_));
dffenr key_r_reg_91_ (.rb(reset), .ck(clk), .d(key_91), .en(n_48), .q(key_r_91_));
dffenr key_r_reg_92_ (.rb(reset), .ck(clk), .d(key_92), .en(n_48), .q(key_r_92_));
dffenr key_r_reg_93_ (.rb(reset), .ck(clk), .d(key_93), .en(n_48), .q(key_r_93_));
dffenr key_r_reg_94_ (.rb(reset), .ck(clk), .d(key_94), .en(n_48), .q(key_r_94_));
dffenr key_r_reg_95_ (.rb(reset), .ck(clk), .d(key_95), .en(n_48), .q(key_r_95_));
dffenr key_r_reg_96_ (.rb(reset), .ck(clk), .d(key_96), .en(n_48), .q(key_r_96_));
dffenr key_r_reg_97_ (.rb(reset), .ck(clk), .d(key_97), .en(n_48), .q(key_r_97_));
dffenr key_r_reg_98_ (.rb(reset), .ck(clk), .d(key_98), .en(n_48), .q(key_r_98_));
dffenr key_r_reg_99_ (.rb(reset), .ck(clk), .d(key_99), .en(n_48), .q(key_r_99_));
dffenr key_r_reg_100_ (.rb(reset), .ck(clk), .d(key_100), .en(n_48), .q(key_r_100_));
dffenr key_r_reg_101_ (.rb(reset), .ck(clk), .d(key_101), .en(n_48), .q(key_r_101_));
dffenr key_r_reg_102_ (.rb(reset), .ck(clk), .d(key_102), .en(n_48), .q(key_r_102_));
dffenr key_r_reg_103_ (.rb(reset), .ck(clk), .d(key_103), .en(n_48), .q(key_r_103_));
dffenr key_r_reg_104_ (.rb(reset), .ck(clk), .d(key_104), .en(n_48), .q(key_r_104_));
dffenr key_r_reg_105_ (.rb(reset), .ck(clk), .d(key_105), .en(n_48), .q(key_r_105_));
dffenr key_r_reg_106_ (.rb(reset), .ck(clk), .d(key_106), .en(n_48), .q(key_r_106_));
dffenr key_r_reg_107_ (.rb(reset), .ck(clk), .d(key_107), .en(n_48), .q(key_r_107_));
dffenr key_r_reg_108_ (.rb(reset), .ck(clk), .d(key_108), .en(n_48), .q(key_r_108_));
dffenr key_r_reg_109_ (.rb(reset), .ck(clk), .d(key_109), .en(n_48), .q(key_r_109_));
dffenr key_r_reg_110_ (.rb(reset), .ck(clk), .d(key_110), .en(n_48), .q(key_r_110_));
dffenr key_r_reg_111_ (.rb(reset), .ck(clk), .d(key_111), .en(n_48), .q(key_r_111_));
dffenr key_r_reg_112_ (.rb(reset), .ck(clk), .d(key_112), .en(n_48), .q(key_r_112_));
dffenr key_r_reg_113_ (.rb(reset), .ck(clk), .d(key_113), .en(n_48), .q(key_r_113_));
dffenr key_r_reg_114_ (.rb(reset), .ck(clk), .d(key_114), .en(n_48), .q(key_r_114_));
dffenr key_r_reg_115_ (.rb(reset), .ck(clk), .d(key_115), .en(n_48), .q(key_r_115_));
dffenr key_r_reg_116_ (.rb(reset), .ck(clk), .d(key_116), .en(n_48), .q(key_r_116_));
dffenr key_r_reg_117_ (.rb(reset), .ck(clk), .d(key_117), .en(n_48), .q(key_r_117_));
dffenr key_r_reg_118_ (.rb(reset), .ck(clk), .d(key_118), .en(n_48), .q(key_r_118_));
dffenr key_r_reg_119_ (.rb(reset), .ck(clk), .d(key_119), .en(n_48), .q(key_r_119_));
dffenr key_r_reg_120_ (.rb(reset), .ck(clk), .d(key_120), .en(n_48), .q(key_r_120_));
dffenr key_r_reg_121_ (.rb(reset), .ck(clk), .d(key_121), .en(n_48), .q(key_r_121_));
dffenr key_r_reg_122_ (.rb(reset), .ck(clk), .d(key_122), .en(n_48), .q(key_r_122_));
dffenr key_r_reg_123_ (.rb(reset), .ck(clk), .d(key_123), .en(n_48), .q(key_r_123_));
dffenr key_r_reg_124_ (.rb(reset), .ck(clk), .d(key_124), .en(n_48), .q(key_r_124_));
dffenr key_r_reg_125_ (.rb(reset), .ck(clk), .d(key_125), .en(n_48), .q(key_r_125_));
dffenr key_r_reg_126_ (.rb(reset), .ck(clk), .d(key_126), .en(n_48), .q(key_r_126_));
dffenr key_r_reg_127_ (.rb(reset), .ck(clk), .d(key_127), .en(n_48), .q(key_r_127_));
dffr ps_reg_0_ (.rb(reset), .ck(clk), .d(n_164), .q(ps_0_));
dffr ps_reg_1_ (.rb(reset), .ck(clk), .d(n_79), .q(ps_1_));
dffr sum_reg_1_ (.rb(reset), .ck(clk), .d(n_78), .q(sum_1_));
dffr sum_reg_2_ (.rb(reset), .ck(clk), .d(n_49), .q(sum_2_));
dffr sum_reg_3_ (.rb(reset), .ck(clk), .d(n_77), .q(sum_3_));
dffr sum_reg_4_ (.rb(reset), .ck(clk), .d(n_76), .q(sum_4_));
dffr sum_reg_5_ (.rb(reset), .ck(clk), .d(n_75), .q(sum_5_));
dffr sum_reg_6_ (.rb(reset), .ck(clk), .d(n_74), .q(sum_6_));
dffr sum_reg_7_ (.rb(reset), .ck(clk), .d(n_73), .q(sum_7_));
dffr sum_reg_8_ (.rb(reset), .ck(clk), .d(n_72), .q(sum_8_));
dffr sum_reg_9_ (.rb(reset), .ck(clk), .d(n_71), .q(sum_9_));
dffr sum_reg_10_ (.rb(reset), .ck(clk), .d(n_50), .q(sum_10_));
dffr sum_reg_11_ (.rb(reset), .ck(clk), .d(n_59), .q(sum_11_));
dffr sum_reg_12_ (.rb(reset), .ck(clk), .d(n_69), .q(sum_12_));
dffr sum_reg_13_ (.rb(reset), .ck(clk), .d(n_68), .q(sum_13_));
dffr sum_reg_14_ (.rb(reset), .ck(clk), .d(n_67), .q(sum_14_));
dffr sum_reg_15_ (.rb(reset), .ck(clk), .d(n_66), .q(sum_15_));
dffr sum_reg_16_ (.rb(reset), .ck(clk), .d(n_65), .q(sum_16_));
dffr sum_reg_17_ (.rb(reset), .ck(clk), .d(n_64), .q(sum_17_));
dffr sum_reg_18_ (.rb(reset), .ck(clk), .d(n_63), .q(sum_18_));
dffr sum_reg_19_ (.rb(reset), .ck(clk), .d(n_62), .q(sum_19_));
dffr sum_reg_20_ (.rb(reset), .ck(clk), .d(n_61), .q(sum_20_));
dffr sum_reg_21_ (.rb(reset), .ck(clk), .d(n_60), .q(sum_21_));
dffr sum_reg_22_ (.rb(reset), .ck(clk), .d(n_70), .q(sum_22_));
dffr sum_reg_23_ (.rb(reset), .ck(clk), .d(n_58), .q(sum_23_));
dffr sum_reg_24_ (.rb(reset), .ck(clk), .d(n_57), .q(sum_24_));
dffr sum_reg_25_ (.rb(reset), .ck(clk), .d(n_56), .q(sum_25_));
dffr sum_reg_26_ (.rb(reset), .ck(clk), .d(n_55), .q(sum_26_));
dffr sum_reg_27_ (.rb(reset), .ck(clk), .d(n_54), .q(sum_27_));
dffr sum_reg_28_ (.rb(reset), .ck(clk), .d(n_53), .q(sum_28_));
dffr sum_reg_29_ (.rb(reset), .ck(clk), .d(n_52), .q(sum_29_));
dffr sum_reg_30_ (.rb(reset), .ck(clk), .d(n_82), .q(sum_30_));
dffr sum_reg_31_ (.rb(reset), .ck(clk), .d(n_51), .q(sum_31_));
dffenr v0_r_reg_0_ (.rb(reset), .ck(clk), .d(in_enc_32), .en(n_48), .q(v0_r_0_));
dffenr v0_r_reg_1_ (.rb(reset), .ck(clk), .d(in_enc_33), .en(n_48), .q(v0_r_1_));
dffenr v0_r_reg_2_ (.rb(reset), .ck(clk), .d(in_enc_34), .en(n_48), .q(v0_r_2_));
dffenr v0_r_reg_3_ (.rb(reset), .ck(clk), .d(in_enc_35), .en(n_48), .q(v0_r_3_));
dffenr v0_r_reg_4_ (.rb(reset), .ck(clk), .d(in_enc_36), .en(n_48), .q(v0_r_4_));
dffenr v0_r_reg_5_ (.rb(reset), .ck(clk), .d(in_enc_37), .en(n_48), .q(v0_r_5_));
dffenr v0_r_reg_6_ (.rb(reset), .ck(clk), .d(in_enc_38), .en(n_48), .q(v0_r_6_));
dffenr v0_r_reg_7_ (.rb(reset), .ck(clk), .d(in_enc_39), .en(n_48), .q(v0_r_7_));
dffenr v0_r_reg_8_ (.rb(reset), .ck(clk), .d(in_enc_40), .en(n_48), .q(v0_r_8_));
dffenr v0_r_reg_9_ (.rb(reset), .ck(clk), .d(in_enc_41), .en(n_48), .q(v0_r_9_));
dffenr v0_r_reg_10_ (.rb(reset), .ck(clk), .d(in_enc_42), .en(n_48), .q(v0_r_10_));
dffenr v0_r_reg_11_ (.rb(reset), .ck(clk), .d(in_enc_43), .en(n_48), .q(v0_r_11_));
dffenr v0_r_reg_12_ (.rb(reset), .ck(clk), .d(in_enc_44), .en(n_48), .q(v0_r_12_));
dffenr v0_r_reg_13_ (.rb(reset), .ck(clk), .d(in_enc_45), .en(n_48), .q(v0_r_13_));
dffenr v0_r_reg_14_ (.rb(reset), .ck(clk), .d(in_enc_46), .en(n_48), .q(v0_r_14_));
dffenr v0_r_reg_15_ (.rb(reset), .ck(clk), .d(in_enc_47), .en(n_48), .q(v0_r_15_));
dffenr v0_r_reg_16_ (.rb(reset), .ck(clk), .d(in_enc_48), .en(n_48), .q(v0_r_16_));
dffenr v0_r_reg_17_ (.rb(reset), .ck(clk), .d(in_enc_49), .en(n_48), .q(v0_r_17_));
dffenr v0_r_reg_18_ (.rb(reset), .ck(clk), .d(in_enc_50), .en(n_48), .q(v0_r_18_));
dffenr v0_r_reg_19_ (.rb(reset), .ck(clk), .d(in_enc_51), .en(n_48), .q(v0_r_19_));
dffenr v0_r_reg_20_ (.rb(reset), .ck(clk), .d(in_enc_52), .en(n_48), .q(v0_r_20_));
dffenr v0_r_reg_21_ (.rb(reset), .ck(clk), .d(in_enc_53), .en(n_48), .q(v0_r_21_));
dffenr v0_r_reg_22_ (.rb(reset), .ck(clk), .d(in_enc_54), .en(n_48), .q(v0_r_22_));
dffenr v0_r_reg_23_ (.rb(reset), .ck(clk), .d(in_enc_55), .en(n_48), .q(v0_r_23_));
dffenr v0_r_reg_24_ (.rb(reset), .ck(clk), .d(in_enc_56), .en(n_48), .q(v0_r_24_));
dffenr v0_r_reg_25_ (.rb(reset), .ck(clk), .d(in_enc_57), .en(n_48), .q(v0_r_25_));
dffenr v0_r_reg_26_ (.rb(reset), .ck(clk), .d(in_enc_58), .en(n_48), .q(v0_r_26_));
dffenr v0_r_reg_27_ (.rb(reset), .ck(clk), .d(in_enc_59), .en(n_48), .q(v0_r_27_));
dffenr v0_r_reg_28_ (.rb(reset), .ck(clk), .d(in_enc_60), .en(n_48), .q(v0_r_28_));
dffenr v0_r_reg_29_ (.rb(reset), .ck(clk), .d(in_enc_61), .en(n_48), .q(v0_r_29_));
dffenr v0_r_reg_30_ (.rb(reset), .ck(clk), .d(in_enc_62), .en(n_48), .q(v0_r_30_));
dffenr v0_r_reg_31_ (.rb(reset), .ck(clk), .d(in_enc_63), .en(n_48), .q(v0_r_31_));
dffr v0_reg_0_ (.rb(reset), .ck(clk), .d(n_163), .q(v0_0_));
dffr v0_reg_1_ (.rb(reset), .ck(clk), .d(n_162), .q(v0_1_));
dffr v0_reg_2_ (.rb(reset), .ck(clk), .d(n_161), .q(v0_2_));
dffr v0_reg_3_ (.rb(reset), .ck(clk), .d(n_160), .q(v0_3_));
dffr v0_reg_4_ (.rb(reset), .ck(clk), .d(n_159), .q(v0_4_));
dffr v0_reg_5_ (.rb(reset), .ck(clk), .d(n_158), .q(v0_5_));
dffr v0_reg_6_ (.rb(reset), .ck(clk), .d(n_157), .q(v0_6_));
dffr v0_reg_7_ (.rb(reset), .ck(clk), .d(n_156), .q(v0_7_));
dffr v0_reg_8_ (.rb(reset), .ck(clk), .d(n_174), .q(v0_8_));
dffr v0_reg_9_ (.rb(reset), .ck(clk), .d(n_175), .q(v0_9_));
dffr v0_reg_10_ (.rb(reset), .ck(clk), .d(n_128), .q(v0_10_));
dffr v0_reg_11_ (.rb(reset), .ck(clk), .d(n_154), .q(v0_11_));
dffr v0_reg_12_ (.rb(reset), .ck(clk), .d(n_153), .q(v0_12_));
dffr v0_reg_13_ (.rb(reset), .ck(clk), .d(n_152), .q(v0_13_));
dffr v0_reg_14_ (.rb(reset), .ck(clk), .d(n_151), .q(v0_14_));
dffr v0_reg_15_ (.rb(reset), .ck(clk), .d(n_150), .q(v0_15_));
dffr v0_reg_16_ (.rb(reset), .ck(clk), .d(n_149), .q(v0_16_));
dffr v0_reg_17_ (.rb(reset), .ck(clk), .d(n_148), .q(v0_17_));
dffr v0_reg_18_ (.rb(reset), .ck(clk), .d(n_147), .q(v0_18_));
dffr v0_reg_19_ (.rb(reset), .ck(clk), .d(n_146), .q(v0_19_));
dffr v0_reg_20_ (.rb(reset), .ck(clk), .d(n_145), .q(v0_20_));
dffr v0_reg_21_ (.rb(reset), .ck(clk), .d(n_144), .q(v0_21_));
dffr v0_reg_22_ (.rb(reset), .ck(clk), .d(n_143), .q(v0_22_));
dffr v0_reg_23_ (.rb(reset), .ck(clk), .d(n_142), .q(v0_23_));
dffr v0_reg_24_ (.rb(reset), .ck(clk), .d(n_141), .q(v0_24_));
dffr v0_reg_25_ (.rb(reset), .ck(clk), .d(n_140), .q(v0_25_));
dffr v0_reg_26_ (.rb(reset), .ck(clk), .d(n_139), .q(v0_26_));
dffr v0_reg_27_ (.rb(reset), .ck(clk), .d(n_138), .q(v0_27_));
dffr v0_reg_28_ (.rb(reset), .ck(clk), .d(n_137), .q(v0_28_));
dffr v0_reg_29_ (.rb(reset), .ck(clk), .d(n_136), .q(v0_29_));
dffr v0_reg_30_ (.rb(reset), .ck(clk), .d(n_135), .q(v0_30_));
dffr v0_reg_31_ (.rb(reset), .ck(clk), .d(n_134), .q(v0_31_));
dffenr v1_r_reg_0_ (.rb(reset), .ck(clk), .d(in_enc_0), .en(n_48), .q(v1_r_0_));
dffenr v1_r_reg_1_ (.rb(reset), .ck(clk), .d(in_enc_1), .en(n_48), .q(v1_r_1_));
dffenr v1_r_reg_2_ (.rb(reset), .ck(clk), .d(in_enc_2), .en(n_48), .q(v1_r_2_));
dffenr v1_r_reg_3_ (.rb(reset), .ck(clk), .d(in_enc_3), .en(n_48), .q(v1_r_3_));
dffenr v1_r_reg_4_ (.rb(reset), .ck(clk), .d(in_enc_4), .en(n_48), .q(v1_r_4_));
dffenr v1_r_reg_5_ (.rb(reset), .ck(clk), .d(in_enc_5), .en(n_48), .q(v1_r_5_));
dffenr v1_r_reg_6_ (.rb(reset), .ck(clk), .d(in_enc_6), .en(n_48), .q(v1_r_6_));
dffenr v1_r_reg_7_ (.rb(reset), .ck(clk), .d(in_enc_7), .en(n_48), .q(v1_r_7_));
dffenr v1_r_reg_8_ (.rb(reset), .ck(clk), .d(in_enc_8), .en(n_48), .q(v1_r_8_));
dffenr v1_r_reg_9_ (.rb(reset), .ck(clk), .d(in_enc_9), .en(n_48), .q(v1_r_9_));
dffenr v1_r_reg_10_ (.rb(reset), .ck(clk), .d(in_enc_10), .en(n_48), .q(v1_r_10_));
dffenr v1_r_reg_11_ (.rb(reset), .ck(clk), .d(in_enc_11), .en(n_48), .q(v1_r_11_));
dffenr v1_r_reg_12_ (.rb(reset), .ck(clk), .d(in_enc_12), .en(n_48), .q(v1_r_12_));
dffenr v1_r_reg_13_ (.rb(reset), .ck(clk), .d(in_enc_13), .en(n_48), .q(v1_r_13_));
dffenr v1_r_reg_14_ (.rb(reset), .ck(clk), .d(in_enc_14), .en(n_48), .q(v1_r_14_));
dffenr v1_r_reg_15_ (.rb(reset), .ck(clk), .d(in_enc_15), .en(n_48), .q(v1_r_15_));
dffenr v1_r_reg_16_ (.rb(reset), .ck(clk), .d(in_enc_16), .en(n_48), .q(v1_r_16_));
dffenr v1_r_reg_17_ (.rb(reset), .ck(clk), .d(in_enc_17), .en(n_48), .q(v1_r_17_));
dffenr v1_r_reg_18_ (.rb(reset), .ck(clk), .d(in_enc_18), .en(n_48), .q(v1_r_18_));
dffenr v1_r_reg_19_ (.rb(reset), .ck(clk), .d(in_enc_19), .en(n_48), .q(v1_r_19_));
dffenr v1_r_reg_20_ (.rb(reset), .ck(clk), .d(in_enc_20), .en(n_48), .q(v1_r_20_));
dffenr v1_r_reg_21_ (.rb(reset), .ck(clk), .d(in_enc_21), .en(n_48), .q(v1_r_21_));
dffenr v1_r_reg_22_ (.rb(reset), .ck(clk), .d(in_enc_22), .en(n_48), .q(v1_r_22_));
dffenr v1_r_reg_23_ (.rb(reset), .ck(clk), .d(in_enc_23), .en(n_48), .q(v1_r_23_));
dffenr v1_r_reg_24_ (.rb(reset), .ck(clk), .d(in_enc_24), .en(n_48), .q(v1_r_24_));
dffenr v1_r_reg_25_ (.rb(reset), .ck(clk), .d(in_enc_25), .en(n_48), .q(v1_r_25_));
dffenr v1_r_reg_26_ (.rb(reset), .ck(clk), .d(in_enc_26), .en(n_48), .q(v1_r_26_));
dffenr v1_r_reg_27_ (.rb(reset), .ck(clk), .d(in_enc_27), .en(n_48), .q(v1_r_27_));
dffenr v1_r_reg_28_ (.rb(reset), .ck(clk), .d(in_enc_28), .en(n_48), .q(v1_r_28_));
dffenr v1_r_reg_29_ (.rb(reset), .ck(clk), .d(in_enc_29), .en(n_48), .q(v1_r_29_));
dffenr v1_r_reg_30_ (.rb(reset), .ck(clk), .d(in_enc_30), .en(n_48), .q(v1_r_30_));
dffenr v1_r_reg_31_ (.rb(reset), .ck(clk), .d(in_enc_31), .en(n_48), .q(v1_r_31_));
dffr v1_reg_0_ (.rb(reset), .ck(clk), .d(n_133), .q(v1_0_));
dffr v1_reg_1_ (.rb(reset), .ck(clk), .d(n_132), .q(v1_1_));
dffr v1_reg_2_ (.rb(reset), .ck(clk), .d(n_131), .q(v1_2_));
dffr v1_reg_3_ (.rb(reset), .ck(clk), .d(n_4337), .q(v1_3_));
dffr v1_reg_4_ (.rb(reset), .ck(clk), .d(n_129), .q(v1_4_));
dffr v1_reg_5_ (.rb(reset), .ck(clk), .d(n_4405), .q(v1_5_));
dffr v1_reg_6_ (.rb(reset), .ck(clk), .d(n_4370), .q(v1_6_));
dffr v1_reg_7_ (.rb(reset), .ck(clk), .d(n_4411), .q(v1_7_));
dffr v1_reg_8_ (.rb(reset), .ck(clk), .d(n_125), .q(v1_8_));
dffr v1_reg_9_ (.rb(reset), .ck(clk), .d(n_3343), .q(v1_9_));
dffr v1_reg_10_ (.rb(reset), .ck(clk), .d(n_3332), .q(v1_10_));
dffr v1_reg_11_ (.rb(reset), .ck(clk), .d(n_3349), .q(v1_11_));
dffr v1_reg_12_ (.rb(reset), .ck(clk), .d(n_3355), .q(v1_12_));
dffr v1_reg_13_ (.rb(reset), .ck(clk), .d(n_4552), .q(v1_13_));
dffr v1_reg_14_ (.rb(reset), .ck(clk), .d(n_3361), .q(v1_14_));
dffr v1_reg_15_ (.rb(reset), .ck(clk), .d(n_3380), .q(v1_15_));
dffr v1_reg_16_ (.rb(reset), .ck(clk), .d(n_117), .q(v1_16_));
dffr v1_reg_17_ (.rb(reset), .ck(clk), .d(n_2391), .q(v1_17_));
dffr v1_reg_18_ (.rb(reset), .ck(clk), .d(n_2406), .q(v1_18_));
dffr v1_reg_19_ (.rb(reset), .ck(clk), .d(n_2421), .q(v1_19_));
dffr v1_reg_20_ (.rb(reset), .ck(clk), .d(n_2433), .q(v1_20_));
dffr v1_reg_21_ (.rb(reset), .ck(clk), .d(n_2448), .q(v1_21_));
dffr v1_reg_22_ (.rb(reset), .ck(clk), .d(n_2463), .q(v1_22_));
dffr v1_reg_23_ (.rb(reset), .ck(clk), .d(n_2478), .q(v1_23_));
dffr v1_reg_24_ (.rb(reset), .ck(clk), .d(n_2493), .q(v1_24_));
dffr v1_reg_25_ (.rb(reset), .ck(clk), .d(n_1731), .q(v1_25_));
dffr v1_reg_26_ (.rb(reset), .ck(clk), .d(n_1756), .q(v1_26_));
dffr v1_reg_27_ (.rb(reset), .ck(clk), .d(n_2498), .q(v1_27_));
dffr v1_reg_28_ (.rb(reset), .ck(clk), .d(n_2506), .q(v1_28_));
dffr v1_reg_29_ (.rb(reset), .ck(clk), .d(n_1691), .q(v1_29_));
dffr v1_reg_30_ (.rb(reset), .ck(clk), .d(n_3625), .q(v1_30_));
dffr v1_reg_31_ (.rb(reset), .ck(clk), .d(n_1710), .q(v1_31_));
mux2 g4167__5703 (.a(v0_r_9_), .b(n_3272), .sel(n_4371), .y(n_175));
mux2 g4189__7114 (.a(v0_r_8_), .b(n_1239), .sel(n_4371), .y(n_174));
nor2 g4190__5266 (.a(n_4371), .b(n_93), .y(n_173));
nor2 g4191__2250 (.a(n_4371), .b(n_101), .y(n_172));
nor2 g4192__6083 (.a(n_99), .b(n_4371), .y(n_171));
nor2 g4194__2703 (.a(n_100), .b(n_4371), .y(n_170));
nor2 g4195__5795 (.a(n_97), .b(n_4371), .y(n_169));
nor2 g4196__7344 (.a(n_98), .b(n_4371), .y(n_168));
nor2 g4197__1840 (.a(n_96), .b(n_4371), .y(n_167));
nor2 g4198__5019 (.a(n_95), .b(n_4371), .y(n_166));
nor2 g4199__1857 (.a(n_94), .b(n_4371), .y(n_165));
nand2 g4200__9906 (.a(n_92), .b(n_47), .y(n_164));
mux2 g4201__8780 (.a(v0_r_0_), .b(n_3269), .sel(n_4371), .y(n_163));
mux2 g4202__4296 (.a(v0_r_1_), .b(n_1246), .sel(n_4371), .y(n_162));
mux2 g4203__3772 (.a(v0_r_2_), .b(n_1245), .sel(n_4371), .y(n_161));
mux2 g4204__1474 (.a(v0_r_3_), .b(n_1244), .sel(n_4371), .y(n_160));
mux2 g4205__4547 (.a(v0_r_4_), .b(n_1243), .sel(n_4371), .y(n_159));
mux2 g4206__9682 (.a(v0_r_5_), .b(n_3139), .sel(n_4371), .y(n_158));
mux2 g4207__2683 (.a(v0_r_6_), .b(n_1241), .sel(n_4371), .y(n_157));
mux2 g4208__1309 (.a(v0_r_7_), .b(n_1240), .sel(n_4371), .y(n_156));
mux2 g4212__2900 (.a(v0_r_11_), .b(n_2005), .sel(n_4371), .y(n_154));
mux2 g4213__2391 (.a(v0_r_12_), .b(n_1235), .sel(n_4371), .y(n_153));
mux2 g4214__7675 (.a(v0_r_13_), .b(n_3580), .sel(n_4371), .y(n_152));
mux2 g4215__7118 (.a(v0_r_14_), .b(n_3708), .sel(n_4371), .y(n_151));
mux2 g4216__8757 (.a(v0_r_15_), .b(n_1998), .sel(n_4371), .y(n_150));
mux2 g4217__1786 (.a(v0_r_16_), .b(n_3713), .sel(n_4371), .y(n_149));
mux2 g4218__5953 (.a(v0_r_17_), .b(n_3490), .sel(n_4371), .y(n_148));
mux2 g4219__5703 (.a(v0_r_18_), .b(n_4048), .sel(n_4371), .y(n_147));
mux2 g4220__7114 (.a(v0_r_19_), .b(n_2195), .sel(n_4371), .y(n_146));
mux2 g4221__5266 (.a(v0_r_20_), .b(n_3687), .sel(n_4371), .y(n_145));
mux2 g4222__2250 (.a(v0_r_21_), .b(n_4306), .sel(n_4371), .y(n_144));
mux2 g4223__6083 (.a(v0_r_22_), .b(n_3505), .sel(n_4371), .y(n_143));
mux2 g4224__2703 (.a(v0_r_23_), .b(n_1224), .sel(n_4371), .y(n_142));
mux2 g4225__5795 (.a(v0_r_24_), .b(n_2033), .sel(n_4371), .y(n_141));
mux2 g4226__7344 (.a(v0_r_25_), .b(n_3611), .sel(n_4371), .y(n_140));
mux2 g4227__1840 (.a(v0_r_26_), .b(n_3502), .sel(n_4371), .y(n_139));
mux2 g4228__5019 (.a(v0_r_27_), .b(n_3525), .sel(n_4371), .y(n_138));
mux2 g4229__1857 (.a(v0_r_28_), .b(n_2586), .sel(n_4371), .y(n_137));
mux2 g4230__9906 (.a(v0_r_29_), .b(n_3914), .sel(n_4371), .y(n_136));
mux2 g4231__8780 (.a(v0_r_30_), .b(n_1217), .sel(n_4371), .y(n_135));
mux2 g4232__4296 (.a(v0_r_31_), .b(n_1216), .sel(n_4371), .y(n_134));
mux2 g4233__3772 (.a(v1_r_0_), .b(n_3144), .sel(n_4371), .y(n_133));
mux2 g4234__1474 (.a(v1_r_1_), .b(n_721), .sel(n_4371), .y(n_132));
mux2 g4235__4547 (.a(v1_r_2_), .b(n_722), .sel(n_4371), .y(n_131));
mux2 g4237__2683 (.a(v1_r_4_), .b(n_724), .sel(n_4371), .y(n_129));
mux2 g4238__1309 (.a(v0_r_10_), .b(n_2961), .sel(n_4371), .y(n_128));
mux2 g4241__2391 (.a(v1_r_8_), .b(n_728), .sel(n_4371), .y(n_125));
mux2 g4249__5266 (.a(v1_r_16_), .b(n_736), .sel(n_4371), .y(n_117));
inv g4265 (.a(n_91), .y(n_101));
inv g4266 (.a(n_90), .y(n_100));
inv g4267 (.a(n_89), .y(n_99));
inv g4269 (.a(n_87), .y(n_98));
inv g4270 (.a(n_86), .y(n_97));
inv g4271 (.a(n_85), .y(n_96));
inv g4272 (.a(n_84), .y(n_95));
inv g4273 (.a(n_83), .y(n_94));
inv g4274 (.a(n_81), .y(n_93));
nand2 g4275__2683 (.a(n_4371), .b(ps_1_), .y(n_92));
nand2 g4276__1309 (.a(n_3112), .b(n_44), .y(n_91));
nand2 g4277__6877 (.a(n_646), .b(n_36), .y(n_90));
nand2 g4278__2900 (.a(n_655), .b(n_38), .y(n_89));
nand2 g4279__2391 (.a(n_652), .b(n_37), .y(n_88));
nand2 g4280__7675 (.a(n_650), .b(n_42), .y(n_87));
nand2 g4281__7118 (.a(n_648), .b(n_39), .y(n_86));
nand2 g4282__8757 (.a(n_654), .b(n_40), .y(n_85));
nand2 g4283__1786 (.a(n_649), .b(n_35), .y(n_84));
nand2 g4284__5953 (.a(n_647), .b(n_45), .y(n_83));
nor2 g4285__5703 (.a(n_30), .b(n_4371), .y(n_82));
nand2 g4286__7114 (.a(n_653), .b(n_46), .y(n_81));
nor2 g4287__5266 (.a(n_4371), .b(sum_0_), .y(n_80));
nand2 g4288__2250 (.a(n_43), .b(n_1800), .y(n_79));
nor2 g4289__6083 (.a(n_4371), .b(n_14), .y(n_78));
nor2 g4290__2703 (.a(n_13), .b(n_4371), .y(n_77));
nor2 g4291__5795 (.a(n_27), .b(n_4371), .y(n_76));
nor2 g4292__7344 (.a(n_31), .b(n_4371), .y(n_75));
nor2 g4293__1840 (.a(n_29), .b(n_4371), .y(n_74));
nor2 g4294__5019 (.a(n_6), .b(n_4371), .y(n_73));
nor2 g4295__1857 (.a(n_7), .b(n_4371), .y(n_72));
nor2 g4296__9906 (.a(n_9), .b(n_4371), .y(n_71));
nor2 g4297__8780 (.a(n_24), .b(n_4371), .y(n_70));
nor2 g4298__4296 (.a(n_3764), .b(n_4371), .y(n_69));
nor2 g4299__3772 (.a(n_21), .b(n_4371), .y(n_68));
nor2 g4300__1474 (.a(n_32), .b(n_4371), .y(n_67));
nor2 g4301__4547 (.a(n_17), .b(n_4371), .y(n_66));
nor2 g4302__9682 (.a(n_8), .b(n_4371), .y(n_65));
nor2 g4303__2683 (.a(n_20), .b(n_4371), .y(n_64));
nor2 g4304__1309 (.a(n_23), .b(n_4371), .y(n_63));
nor2 g4305__6877 (.a(n_3), .b(n_4371), .y(n_62));
nor2 g4306__2900 (.a(n_19), .b(n_4371), .y(n_61));
nor2 g4307__2391 (.a(n_4), .b(n_4371), .y(n_60));
nor2 g4308__7675 (.a(n_3840), .b(n_4371), .y(n_59));
nor2 g4309__7118 (.a(n_26), .b(n_4371), .y(n_58));
nor2 g4310__8757 (.a(n_33), .b(n_4371), .y(n_57));
nor2 g4311__1786 (.a(n_28), .b(n_4371), .y(n_56));
nor2 g4312__5953 (.a(n_16), .b(n_4371), .y(n_55));
nor2 g4313__5703 (.a(n_15), .b(n_4371), .y(n_54));
nor2 g4314__7114 (.a(n_18), .b(n_4371), .y(n_53));
nor2 g4315__5266 (.a(n_5), .b(n_4371), .y(n_52));
nor2 g4316__2250 (.a(n_12), .b(n_4371), .y(n_51));
nor2 g4317__6083 (.a(n_25), .b(n_4371), .y(n_50));
nor2 g4318__2703 (.a(n_4371), .b(n_11), .y(n_49));
inv g4319 (.a(n_48), .y(n_47));
nand2 g4320__5795 (.a(sum_0_), .b(counter_1_), .y(n_46));
nand2 g4321__7344 (.a(n_649), .b(counter_10_), .y(n_45));
nand2 g4322__1840 (.a(n_653), .b(counter_2_), .y(n_44));
nand2 g4323__5019 (.a(n_647), .b(ps_1_), .y(n_43));
nand2 g4324__1857 (.a(n_652), .b(counter_6_), .y(n_42));
nor2 g4325__9906 (.a(ps_0_), .b(ps_1_), .y(n_48));
nand2 g4327__8780 (.a(n_648), .b(counter_8_), .y(n_40));
nand2 g4328__4296 (.a(n_650), .b(counter_7_), .y(n_39));
nand2 g4329__3772 (.a(n_646), .b(counter_4_), .y(n_38));
nand2 g4330__1474 (.a(n_655), .b(counter_5_), .y(n_37));
nand2 g4331__4547 (.a(n_3112), .b(counter_3_), .y(n_36));
nand2 g4332__9682 (.a(n_654), .b(counter_9_), .y(n_35));
inv g4335 (.a(n_1287), .y(n_33));
inv g4336 (.a(n_1297), .y(n_32));
inv g4337 (.a(n_1306), .y(n_31));
inv g4338 (.a(n_1281), .y(n_30));
inv g4339 (.a(n_1305), .y(n_29));
inv g4340 (.a(n_1286), .y(n_28));
inv g4341 (.a(n_1307), .y(n_27));
inv g4342 (.a(n_1288), .y(n_26));
inv g4343 (.a(n_1301), .y(n_25));
inv g4344 (.a(n_1289), .y(n_24));
inv g4345 (.a(n_1293), .y(n_23));
inv g4347 (.a(n_1298), .y(n_21));
inv g4348 (.a(n_1294), .y(n_20));
inv g4349 (.a(n_1291), .y(n_19));
inv g4350 (.a(n_1283), .y(n_18));
inv g4351 (.a(n_1296), .y(n_17));
inv g4352 (.a(n_1285), .y(n_16));
inv g4353 (.a(n_1284), .y(n_15));
inv g4354 (.a(n_2066), .y(n_14));
inv g4355 (.a(n_1308), .y(n_13));
inv g4356 (.a(n_1280), .y(n_12));
inv g4357 (.a(n_2070), .y(n_11));
inv g4359 (.a(n_1302), .y(n_9));
inv g4360 (.a(n_1295), .y(n_8));
inv g4361 (.a(n_1303), .y(n_7));
inv g4362 (.a(n_1304), .y(n_6));
inv g4363 (.a(n_1282), .y(n_5));
inv g4364 (.a(n_1290), .y(n_4));
inv g4365 (.a(n_1292), .y(n_3));
inv g3 (.a(n_1), .y(n_0));
nor2 g2__1309 (.a(n_88), .b(n_4371), .y(n_1));
xor2 g6391__7118 (.a(n_799), .b(n_798), .y(n_797));
xor2 g6394__5953 (.a(n_766), .b(n_765), .y(n_764));
xor2 g6399__6083 (.a(n_942), .b(n_943), .y(n_941));
xor2 g6400__2703 (.a(n_939), .b(n_940), .y(n_938));
xor2 g6428__2703 (.a(n_849), .b(n_850), .y(n_848));
xor2 g6434__9906 (.a(n_796), .b(n_795), .y(n_794));
xor2 g6436__4296 (.a(n_790), .b(n_789), .y(n_788));
xor2 g6439__4547 (.a(n_778), .b(n_777), .y(n_776));
nand2 add_88_69_g1547__2391 (.a(n_3599), .b(add_88_69_n_1270), .y(add_88_69_n_1243));
xor2 add_88_69_g1551__1786 (.a(add_88_69_n_1278), .b(add_88_69_n_1614), .y(n_796));
xor2 add_88_69_g1556__2250 (.a(add_88_69_n_1284), .b(add_88_69_n_1608), .y(n_799));
xor2 add_88_69_g1557__6083 (.a(add_88_69_n_1277), .b(add_88_69_n_1606), .y(n_790));
nand2 add_88_69_g1563__1857 (.a(n_2103), .b(add_88_69_n_1376), .y(add_88_69_n_1259));
nand2 add_88_69_g1564__9906 (.a(n_2103), .b(add_88_69_n_1528), .y(add_88_69_n_1261));
nor2 add_88_69_g1565__8780 (.a(add_88_69_n_1280), .b(add_88_69_n_1378), .y(add_88_69_n_1262));
nor2 add_88_69_g1566__4296 (.a(add_88_69_n_1277), .b(add_88_69_n_1417), .y(add_88_69_n_1263));
nor2 add_88_69_g1567__3772 (.a(add_88_69_n_1280), .b(add_88_69_n_1373), .y(add_88_69_n_1265));
nand2 add_88_69_g1568__1474 (.a(n_2103), .b(add_88_69_n_1398), .y(add_88_69_n_1267));
nand2 add_88_69_g1569__4547 (.a(n_2103), .b(add_88_69_n_1414), .y(add_88_69_n_1268));
nand2 add_88_69_g1571__2683 (.a(n_2103), .b(add_88_69_n_1407), .y(add_88_69_n_1270));
nor2 add_88_69_g1572__1309 (.a(add_88_69_n_1280), .b(add_88_69_n_1422), .y(add_88_69_n_1271));
nor2 add_88_69_g1573__6877 (.a(add_88_69_n_1280), .b(add_88_69_n_1476), .y(add_88_69_n_1272));
nand2 add_88_69_g1575__2391 (.a(n_2103), .b(add_88_69_n_1400), .y(add_88_69_n_1274));
nand2 add_88_69_g1577__7118 (.a(n_2103), .b(add_88_69_n_1508), .y(add_88_69_n_1276));
nor2 add_88_69_g1578__8757 (.a(add_88_69_n_1370), .b(add_88_69_n_1303), .y(add_88_69_n_1277));
nor2 add_88_69_g1579__1786 (.a(add_88_69_n_1321), .b(add_88_69_n_1300), .y(add_88_69_n_1278));
inv add_88_69_g1580 (.a(n_2103), .y(add_88_69_n_1280));
nor2 add_88_69_g1585__2250 (.a(add_88_69_n_1337), .b(add_88_69_n_1302), .y(add_88_69_n_1284));
xor2 add_88_69_g1587__2703 (.a(add_88_69_n_1308), .b(add_88_69_n_1605), .y(n_778));
inv add_88_69_g1589 (.a(add_88_69_n_1293), .y(add_88_69_n_1288));
nor2 add_88_69_g1590__7344 (.a(add_88_69_n_1329), .b(add_88_69_n_1316), .y(add_88_69_n_1289));
nor2 add_88_69_g1591__1840 (.a(add_88_69_n_1334), .b(add_88_69_n_1313), .y(add_88_69_n_1290));
nand2 add_88_69_g1593__1857 (.a(add_88_69_n_1425), .b(add_88_69_n_1309), .y(add_88_69_n_1292));
nor2 add_88_69_g1594__9906 (.a(add_88_69_n_1308), .b(add_88_69_n_1722), .y(add_88_69_n_1293));
nand2 add_88_69_g1595__8780 (.a(add_88_69_n_1309), .b(add_88_69_n_1419), .y(add_88_69_n_1295));
nand2 add_88_69_g1596__4296 (.a(add_88_69_n_1309), .b(add_88_69_n_1525), .y(add_88_69_n_1297));
nand2 add_88_69_g1597__3772 (.a(n_2038), .b(add_88_69_n_1311), .y(add_88_69_n_1298));
nor2 add_88_69_g1599__4547 (.a(add_88_69_n_1447), .b(add_88_69_n_1308), .y(add_88_69_n_1300));
nor2 add_88_69_g1601__2683 (.a(add_88_69_n_1458), .b(add_88_69_n_1308), .y(add_88_69_n_1302));
nor2 add_88_69_g1602__1309 (.a(add_88_69_n_1308), .b(add_88_69_n_1473), .y(add_88_69_n_1303));
nor2 add_88_69_g1603__6877 (.a(add_88_69_n_1308), .b(add_88_69_n_1506), .y(add_88_69_n_1304));
inv add_88_69_g1607 (.a(add_88_69_n_1308), .y(add_88_69_n_1309));
nor2 add_88_69_g1608__7118 (.a(add_88_69_n_1381), .b(add_88_69_n_1330), .y(add_88_69_n_1308));
nand2 add_88_69_g1610__1786 (.a(n_3600), .b(add_88_69_n_1406), .y(add_88_69_n_1311));
nor2 add_88_69_g1611__5953 (.a(n_3599), .b(add_88_69_n_1405), .y(add_88_69_n_1313));
nor2 add_88_69_g1612__5703 (.a(n_3599), .b(add_88_69_n_1477), .y(add_88_69_n_1315));
nor2 add_88_69_g1613__7114 (.a(n_3599), .b(add_88_69_n_1438), .y(add_88_69_n_1316));
nand2 add_88_69_g1615__2250 (.a(n_3901), .b(n_3962), .y(add_88_69_n_1318));
nand2 add_88_69_g1617__6083 (.a(add_88_69_n_1345), .b(add_88_69_n_1499), .y(add_88_69_n_1321));
nor2 add_88_69_g1618__2703 (.a(add_88_69_n_1385), .b(add_88_69_n_1343), .y(add_88_69_n_1322));
nand2 add_88_69_g1619__5795 (.a(add_88_69_n_1515), .b(add_88_69_n_1359), .y(add_88_69_n_1323));
nor2 add_88_69_g1622__5019 (.a(add_88_69_n_1344), .b(add_88_69_n_1638), .y(add_88_69_n_1327));
nand2 add_88_69_g1623__1857 (.a(add_88_69_n_1360), .b(n_4303), .y(add_88_69_n_1328));
nand2 add_88_69_g1624__9906 (.a(add_88_69_n_1358), .b(add_88_69_n_1389), .y(add_88_69_n_1329));
nor2 add_88_69_g1626__4296 (.a(add_88_69_n_1342), .b(add_88_69_n_1518), .y(add_88_69_n_1330));
nor2 add_88_69_g1627__3772 (.a(add_88_69_n_1356), .b(add_88_69_n_1662), .y(add_88_69_n_1331));
xor2 add_88_69_g1629__4547 (.a(add_88_69_n_1601), .b(add_88_69_n_1369), .y(n_766));
nand2 add_88_69_g1630__9682 (.a(add_88_69_n_1347), .b(add_88_69_n_1466), .y(add_88_69_n_1334));
nand2 add_88_69_g1633__6877 (.a(add_88_69_n_1382), .b(add_88_69_n_1364), .y(add_88_69_n_1337));
nor2 add_88_69_g1636__7675 (.a(add_88_69_n_1371), .b(add_88_69_n_1470), .y(add_88_69_n_1343));
nor2 add_88_69_g1637__7118 (.a(add_88_69_n_1367), .b(n_3619), .y(add_88_69_n_1344));
nand2 add_88_69_g1638__8757 (.a(add_88_69_n_1370), .b(add_88_69_n_1531), .y(add_88_69_n_1345));
nand2 add_88_69_g1639__1786 (.a(n_1919), .b(add_88_69_n_1524), .y(add_88_69_n_1347));
nand2 add_88_69_g1642__7114 (.a(add_88_69_n_1366), .b(add_88_69_n_1529), .y(add_88_69_n_1341));
nand2 add_88_69_g1643__5266 (.a(add_88_69_n_1515), .b(add_88_69_n_1369), .y(add_88_69_n_1342));
nand2 add_88_69_g1644__2250 (.a(add_88_69_n_1732), .b(add_88_69_n_1369), .y(add_88_69_n_1355));
nor2 add_88_69_g1645__6083 (.a(add_88_69_n_1371), .b(add_88_69_n_1737), .y(add_88_69_n_1356));
nand2 add_88_69_g1646__2703 (.a(n_1919), .b(add_88_69_n_1492), .y(add_88_69_n_1358));
nor2 add_88_69_g1647__5795 (.a(add_88_69_n_1674), .b(add_88_69_n_1368), .y(add_88_69_n_1359));
nand2 add_88_69_g1648__7344 (.a(add_88_69_n_1385), .b(add_88_69_n_1671), .y(add_88_69_n_1360));
nor2 add_88_69_g1650__5019 (.a(add_88_69_n_1367), .b(add_88_69_n_1464), .y(add_88_69_n_1363));
nand2 add_88_69_g1651__1857 (.a(add_88_69_n_1370), .b(add_88_69_n_1490), .y(add_88_69_n_1364));
inv add_88_69_g1653 (.a(add_88_69_n_1366), .y(add_88_69_n_1367));
inv add_88_69_g1654 (.a(add_88_69_n_1369), .y(add_88_69_n_1368));
inv add_88_69_g1655 (.a(add_88_69_n_1370), .y(add_88_69_n_1371));
nand2 add_88_69_g1656__9906 (.a(add_88_69_n_1439), .b(add_88_69_n_1643), .y(add_88_69_n_1372));
nand2 add_88_69_g1657__8780 (.a(add_88_69_n_1406), .b(add_88_69_n_1407), .y(add_88_69_n_1373));
nor2 add_88_69_g1658__4296 (.a(add_88_69_n_1408), .b(add_88_69_n_1739), .y(add_88_69_n_1376));
nand2 add_88_69_g1659__3772 (.a(add_88_69_n_1404), .b(n_3574), .y(add_88_69_n_1377));
nand2 add_88_69_g1660__1474 (.a(add_88_69_n_1407), .b(add_88_69_n_1530), .y(add_88_69_n_1378));
nor2 add_88_69_g1661__4547 (.a(add_88_69_n_1441), .b(add_88_69_n_1659), .y(add_88_69_n_1380));
nand2 add_88_69_g1662__9682 (.a(add_88_69_n_1443), .b(add_88_69_n_1505), .y(add_88_69_n_1381));
nor2 add_88_69_g1663__2683 (.a(add_88_69_n_1445), .b(add_88_69_n_1734), .y(add_88_69_n_1382));
nand2 add_88_69_g1665__6877 (.a(add_88_69_n_1444), .b(add_88_69_n_1504), .y(add_88_69_n_1366));
nand2 add_88_69_g1666__2900 (.a(add_88_69_n_1479), .b(add_88_69_n_1449), .y(add_88_69_n_1369));
nand2 add_88_69_g1667__2391 (.a(add_88_69_n_1431), .b(add_88_69_n_1481), .y(add_88_69_n_1370));
nor2 add_88_69_g1670__7118 (.a(add_88_69_n_1412), .b(add_88_69_n_1697), .y(add_88_69_n_1389));
nor2 add_88_69_g1674__5703 (.a(add_88_69_n_1408), .b(add_88_69_n_1477), .y(add_88_69_n_1395));
nor2 add_88_69_g1675__7114 (.a(add_88_69_n_1409), .b(add_88_69_n_1654), .y(add_88_69_n_1397));
nor2 add_88_69_g1676__5266 (.a(add_88_69_n_1438), .b(add_88_69_n_1408), .y(add_88_69_n_1398));
nor2 add_88_69_g1677__2250 (.a(add_88_69_n_1405), .b(add_88_69_n_1408), .y(add_88_69_n_1400));
nand2 add_88_69_g1679__2703 (.a(add_88_69_n_1453), .b(add_88_69_n_1510), .y(add_88_69_n_1385));
inv add_88_69_g1682 (.a(n_2843), .y(add_88_69_n_1404));
inv add_88_69_g1683 (.a(add_88_69_n_1407), .y(add_88_69_n_1408));
nor2 add_88_69_g1684__7344 (.a(add_88_69_n_1501), .b(add_88_69_n_1674), .y(add_88_69_n_1409));
nor2 add_88_69_g1685__1840 (.a(add_88_69_n_1466), .b(add_88_69_n_1649), .y(add_88_69_n_1412));
nor2 add_88_69_g1686__5019 (.a(n_3619), .b(add_88_69_n_1476), .y(add_88_69_n_1414));
nand2 add_88_69_g1687__1857 (.a(add_88_69_n_1469), .b(add_88_69_n_1671), .y(add_88_69_n_1417));
nor2 add_88_69_g1688__9906 (.a(add_88_69_n_1473), .b(add_88_69_n_1737), .y(add_88_69_n_1419));
nand2 add_88_69_g1689__8780 (.a(add_88_69_n_1529), .b(add_88_69_n_1475), .y(add_88_69_n_1422));
nand2 add_88_69_g1690__4296 (.a(n_2211), .b(n_2842), .y(add_88_69_n_1424));
nor2 add_88_69_g1691__3772 (.a(add_88_69_n_1470), .b(add_88_69_n_1473), .y(add_88_69_n_1425));
nand2 add_88_69_g1694__9682 (.a(add_88_69_n_1472), .b(add_88_69_n_1516), .y(add_88_69_n_1431));
nand2 add_88_69_g1696__1309 (.a(add_88_69_n_1478), .b(add_88_69_n_1524), .y(add_88_69_n_1405));
nor2 add_88_69_g1697__6877 (.a(add_88_69_n_1477), .b(n_1904), .y(add_88_69_n_1406));
nor2 add_88_69_g1698__2900 (.a(add_88_69_n_1465), .b(add_88_69_n_1476), .y(add_88_69_n_1407));
inv add_88_69_g1699 (.a(add_88_69_n_1454), .y(add_88_69_n_1437));
nand2 add_88_69_g1700__2391 (.a(add_88_69_n_1472), .b(add_88_69_n_1673), .y(add_88_69_n_1439));
nor2 add_88_69_g1701__7675 (.a(n_3887), .b(add_88_69_n_1740), .y(add_88_69_n_1441));
nand2 add_88_69_g1702__7118 (.a(add_88_69_n_1502), .b(add_88_69_n_1519), .y(add_88_69_n_1443));
nand2 add_88_69_g1703__8757 (.a(add_88_69_n_1496), .b(add_88_69_n_1522), .y(add_88_69_n_1444));
nor2 add_88_69_g1704__1786 (.a(add_88_69_n_1499), .b(add_88_69_n_1676), .y(add_88_69_n_1445));
nand2 add_88_69_g1705__5953 (.a(add_88_69_n_1531), .b(add_88_69_n_1474), .y(add_88_69_n_1447));
nand2 add_88_69_g1706__5703 (.a(add_88_69_n_1538), .b(n_3164), .y(add_88_69_n_1449));
nand2 add_88_69_g1708__5266 (.a(n_3164), .b(add_88_69_n_1730), .y(add_88_69_n_1452));
nand2 add_88_69_g1709__2250 (.a(add_88_69_n_1500), .b(add_88_69_n_1520), .y(add_88_69_n_1453));
nor2 add_88_69_g1710__6083 (.a(n_2025), .b(add_88_69_n_1668), .y(add_88_69_n_1454));
nor2 add_88_69_g1711__2703 (.a(add_88_69_n_1464), .b(add_88_69_n_1476), .y(add_88_69_n_1456));
nand2 add_88_69_g1712__5795 (.a(add_88_69_n_1490), .b(add_88_69_n_1474), .y(add_88_69_n_1458));
nand2 add_88_69_g1714__1840 (.a(add_88_69_n_1478), .b(add_88_69_n_1492), .y(add_88_69_n_1438));
inv add_88_69_g1716 (.a(add_88_69_n_1470), .y(add_88_69_n_1469));
inv add_88_69_g1717 (.a(add_88_69_n_1472), .y(add_88_69_n_1471));
inv add_88_69_g1718 (.a(add_88_69_n_1473), .y(add_88_69_n_1474));
inv add_88_69_g1719 (.a(add_88_69_n_1476), .y(add_88_69_n_1475));
inv add_88_69_g1720 (.a(add_88_69_n_1477), .y(add_88_69_n_1478));
nor2 add_88_69_g1721__5019 (.a(add_88_69_n_1548), .b(add_88_69_n_1698), .y(add_88_69_n_1479));
nor2 add_88_69_g1723__9906 (.a(add_88_69_n_1557), .b(add_88_69_n_1708), .y(add_88_69_n_1481));
nand2 add_88_69_g1725__4296 (.a(add_88_69_n_1529), .b(n_2841), .y(add_88_69_n_1464));
nand2 add_88_69_g1726__3772 (.a(n_2842), .b(add_88_69_n_1529), .y(add_88_69_n_1465));
nor2 add_88_69_g1727__1474 (.a(add_88_69_n_1547), .b(add_88_69_n_1704), .y(add_88_69_n_1466));
nand2 add_88_69_g1729__9682 (.a(add_88_69_n_1520), .b(add_88_69_n_1531), .y(add_88_69_n_1470));
nand2 add_88_69_g1730__2683 (.a(add_88_69_n_1513), .b(add_88_69_n_1702), .y(add_88_69_n_1472));
nand2 add_88_69_g1731__1309 (.a(add_88_69_n_1516), .b(add_88_69_n_1525), .y(add_88_69_n_1473));
nand2 add_88_69_g1732__6877 (.a(add_88_69_n_1522), .b(add_88_69_n_1528), .y(add_88_69_n_1476));
nand2 add_88_69_g1733__2900 (.a(add_88_69_n_1530), .b(n_1917), .y(add_88_69_n_1477));
inv add_88_69_g1735 (.a(n_3887), .y(add_88_69_n_1496));
inv add_88_69_g1737 (.a(add_88_69_n_1499), .y(add_88_69_n_1500));
inv add_88_69_g1738 (.a(add_88_69_n_1501), .y(add_88_69_n_1502));
nor2 add_88_69_g1739__2391 (.a(add_88_69_n_1551), .b(add_88_69_n_1631), .y(add_88_69_n_1504));
nor2 add_88_69_g1740__7675 (.a(add_88_69_n_1543), .b(add_88_69_n_1711), .y(add_88_69_n_1505));
nand2 add_88_69_g1741__7118 (.a(add_88_69_n_1525), .b(add_88_69_n_1673), .y(add_88_69_n_1506));
nor2 add_88_69_g1742__8757 (.a(add_88_69_n_1527), .b(add_88_69_n_1740), .y(add_88_69_n_1508));
nor2 add_88_69_g1743__1786 (.a(add_88_69_n_1556), .b(add_88_69_n_1706), .y(add_88_69_n_1510));
nor2 add_88_69_g1744__5953 (.a(add_88_69_n_1532), .b(add_88_69_n_1676), .y(add_88_69_n_1490));
nand2 add_88_69_g1745__5703 (.a(add_88_69_n_1530), .b(add_88_69_n_1669), .y(add_88_69_n_1491));
nor2 add_88_69_g1746__7114 (.a(add_88_69_n_1523), .b(add_88_69_n_1649), .y(add_88_69_n_1492));
nor2 add_88_69_g1750__2703 (.a(add_88_69_n_1535), .b(add_88_69_n_1710), .y(add_88_69_n_1499));
nor2 add_88_69_g1751__5795 (.a(add_88_69_n_1545), .b(add_88_69_n_1700), .y(add_88_69_n_1501));
inv add_88_69_g1753 (.a(add_88_69_n_1536), .y(add_88_69_n_1513));
inv add_88_69_g1754 (.a(add_88_69_n_1554), .y(add_88_69_n_1514));
inv add_88_69_g1755 (.a(add_88_69_n_1519), .y(add_88_69_n_1518));
inv add_88_69_g1756 (.a(add_88_69_n_1524), .y(add_88_69_n_1523));
inv add_88_69_g1757 (.a(add_88_69_n_1528), .y(add_88_69_n_1527));
inv add_88_69_g1758 (.a(add_88_69_n_1531), .y(add_88_69_n_1532));
nor2 add_88_69_g1760__5019 (.a(add_88_69_n_1663), .b(n_2730), .y(add_88_69_n_1535));
nor2 add_88_69_g1761__1857 (.a(add_88_69_n_1723), .b(add_88_69_n_1714), .y(add_88_69_n_1536));
nor2 add_88_69_g1762__9906 (.a(add_88_69_n_1718), .b(add_88_69_n_1729), .y(add_88_69_n_1538));
nor2 add_88_69_g1765__3772 (.a(add_88_69_n_1655), .b(add_88_69_n_1653), .y(add_88_69_n_1543));
nor2 add_88_69_g1767__4547 (.a(add_88_69_n_1728), .b(add_88_69_n_1646), .y(add_88_69_n_1545));
nor2 add_88_69_g1768__9682 (.a(n_2034), .b(add_88_69_n_1716), .y(add_88_69_n_1547));
nor2 add_88_69_g1769__2683 (.a(add_88_69_n_1644), .b(add_88_69_n_1718), .y(add_88_69_n_1548));
nor2 add_88_69_g1770__1309 (.a(add_88_69_n_1660), .b(add_88_69_n_1650), .y(add_88_69_n_1551));
nor2 add_88_69_g1772__2900 (.a(n_3157), .b(add_88_69_n_1636), .y(add_88_69_n_1554));
nor2 add_88_69_g1773__2391 (.a(add_88_69_n_1735), .b(n_3444), .y(add_88_69_n_1556));
nor2 add_88_69_g1774__7675 (.a(add_88_69_n_1643), .b(add_88_69_n_1720), .y(add_88_69_n_1557));
nor2 add_88_69_g1775__7118 (.a(add_88_69_n_1646), .b(add_88_69_n_1731), .y(add_88_69_n_1515));
nor2 add_88_69_g1776__8757 (.a(add_88_69_n_1672), .b(add_88_69_n_1720), .y(add_88_69_n_1516));
nor2 add_88_69_g1779__5703 (.a(add_88_69_n_1653), .b(add_88_69_n_1674), .y(add_88_69_n_1519));
nor2 add_88_69_g1780__7114 (.a(n_3444), .b(add_88_69_n_1676), .y(add_88_69_n_1520));
nor2 add_88_69_g1782__2250 (.a(add_88_69_n_1650), .b(add_88_69_n_1740), .y(add_88_69_n_1522));
nor2 add_88_69_g1783 (.a(add_88_69_n_1716), .b(n_1904), .y(add_88_69_n_1524));
nor2 add_88_69_g1784 (.a(add_88_69_n_1714), .b(add_88_69_n_1722), .y(add_88_69_n_1525));
nor2 add_88_69_g1786 (.a(n_3454), .b(add_88_69_n_1670), .y(add_88_69_n_1528));
nor2 add_88_69_g1787 (.a(n_2096), .b(n_3619), .y(add_88_69_n_1529));
nor2 add_88_69_g1788 (.a(add_88_69_n_1647), .b(add_88_69_n_1739), .y(add_88_69_n_1530));
nor2 add_88_69_g1789 (.a(n_2730), .b(add_88_69_n_1737), .y(add_88_69_n_1531));
nor2 add_88_69_g1803 (.a(add_88_69_n_1727), .b(add_88_69_n_1731), .y(add_88_69_n_1601));
nand2 add_88_69_g1806 (.a(add_88_69_n_1723), .b(add_88_69_n_1721), .y(add_88_69_n_1605));
nand2 add_88_69_g1807 (.a(add_88_69_n_1663), .b(add_88_69_n_1736), .y(add_88_69_n_1606));
nand2 add_88_69_g1808 (.a(n_4090), .b(add_88_69_n_1725), .y(add_88_69_n_1608));
nor2 add_88_69_g1811 (.a(add_88_69_n_1712), .b(add_88_69_n_1670), .y(add_88_69_n_1612));
nand2 add_88_69_g1812 (.a(add_88_69_n_1735), .b(add_88_69_n_1675), .y(add_88_69_n_1614));
inv add_88_69_g1822 (.a(add_88_69_n_1679), .y(add_88_69_n_1631));
inv add_88_69_g1823 (.a(add_88_69_n_1633), .y(add_88_69_n_1632));
inv add_88_69_g1824 (.a(add_88_69_n_1680), .y(add_88_69_n_1634));
inv add_88_69_g1825 (.a(add_88_69_n_1636), .y(add_88_69_n_1635));
inv add_88_69_g1826 (.a(n_2520), .y(add_88_69_n_1638));
inv add_88_69_g1828 (.a(add_88_69_n_1643), .y(add_88_69_n_1642));
inv add_88_69_g1829 (.a(add_88_69_n_1644), .y(add_88_69_n_1645));
inv add_88_69_g1831 (.a(add_88_69_n_1655), .y(add_88_69_n_1654));
inv add_88_69_g1832 (.a(n_3454), .y(add_88_69_n_1656));
inv add_88_69_g1833 (.a(add_88_69_n_1660), .y(add_88_69_n_1659));
inv add_88_69_g1834 (.a(add_88_69_n_1663), .y(add_88_69_n_1662));
inv add_88_69_g1837 (.a(add_88_69_n_1668), .y(add_88_69_n_1669));
inv add_88_69_g1838 (.a(add_88_69_n_1670), .y(add_88_69_n_1671));
inv add_88_69_g1839 (.a(add_88_69_n_1672), .y(add_88_69_n_1673));
inv add_88_69_g1840 (.a(add_88_69_n_1676), .y(add_88_69_n_1675));
nand2 add_88_69_g1842 (.a(n_974), .b(n_2195), .y(add_88_69_n_1679));
nand2 add_88_69_g1843 (.a(n_2610), .b(n_3490), .y(add_88_69_n_1633));
nand2 add_88_69_g1844 (.a(n_2588), .b(n_1224), .y(add_88_69_n_1680));
nor2 add_88_69_g1845 (.a(n_1241), .b(n_1246), .y(add_88_69_n_1636));
nand2 add_88_69_g1849 (.a(n_983), .b(n_2961), .y(add_88_69_n_1643));
nand2 add_88_69_g1850 (.a(n_1240), .b(n_1245), .y(add_88_69_n_1644));
nor2 add_88_69_g1851 (.a(n_988), .b(n_3139), .y(add_88_69_n_1646));
nor2 add_88_69_g1852 (.a(n_968), .b(n_3611), .y(add_88_69_n_1647));
nor2 add_88_69_g1853 (.a(n_3525), .b(n_1224), .y(add_88_69_n_1648));
nor2 add_88_69_g1854 (.a(n_1217), .b(n_3502), .y(add_88_69_n_1649));
nor2 add_88_69_g1855 (.a(n_974), .b(n_2195), .y(add_88_69_n_1650));
nor2 add_88_69_g1857 (.a(n_986), .b(n_1240), .y(add_88_69_n_1653));
nand2 add_88_69_g1858 (.a(n_987), .b(n_1241), .y(add_88_69_n_1655));
nand2 add_88_69_g1861 (.a(n_975), .b(n_4048), .y(add_88_69_n_1660));
nand2 add_88_69_g1863 (.a(n_981), .b(n_1235), .y(add_88_69_n_1663));
nor2 add_88_69_g1866 (.a(n_967), .b(n_3502), .y(add_88_69_n_1668));
nor2 add_88_69_g1867 (.a(n_3888), .b(n_3713), .y(add_88_69_n_1670));
nor2 add_88_69_g1868 (.a(n_983), .b(n_2961), .y(add_88_69_n_1672));
nor2 add_88_69_g1869 (.a(n_987), .b(n_1241), .y(add_88_69_n_1674));
nor2 add_88_69_g1870 (.a(n_2194), .b(n_3708), .y(add_88_69_n_1676));
inv add_88_69_g1871 (.a(add_88_69_n_1743), .y(add_88_69_n_1697));
inv add_88_69_g1872 (.a(add_88_69_n_1745), .y(add_88_69_n_1698));
inv add_88_69_g1873 (.a(add_88_69_n_1746), .y(add_88_69_n_1699));
inv add_88_69_g1874 (.a(add_88_69_n_1749), .y(add_88_69_n_1700));
inv add_88_69_g1875 (.a(add_88_69_n_1702), .y(add_88_69_n_1701));
inv add_88_69_g1876 (.a(add_88_69_n_1705), .y(add_88_69_n_1704));
inv add_88_69_g1877 (.a(n_4090), .y(add_88_69_n_1706));
inv add_88_69_g1878 (.a(add_88_69_n_1709), .y(add_88_69_n_1708));
inv add_88_69_g1879 (.a(add_88_69_n_1752), .y(add_88_69_n_1710));
inv add_88_69_g1880 (.a(add_88_69_n_1755), .y(add_88_69_n_1711));
inv add_88_69_g1881 (.a(n_4303), .y(add_88_69_n_1712));
inv add_88_69_g1882 (.a(add_88_69_n_1716), .y(add_88_69_n_1715));
inv add_88_69_g1883 (.a(add_88_69_n_1720), .y(add_88_69_n_1719));
inv add_88_69_g1884 (.a(add_88_69_n_1722), .y(add_88_69_n_1721));
inv add_88_69_g1885 (.a(n_3444), .y(add_88_69_n_1725));
inv add_88_69_g1886 (.a(add_88_69_n_1728), .y(add_88_69_n_1727));
inv add_88_69_g1887 (.a(add_88_69_n_1729), .y(add_88_69_n_1730));
inv add_88_69_g1888 (.a(add_88_69_n_1731), .y(add_88_69_n_1732));
inv add_88_69_g1889 (.a(add_88_69_n_1735), .y(add_88_69_n_1734));
inv add_88_69_g1890 (.a(add_88_69_n_1737), .y(add_88_69_n_1736));
inv add_88_69_g1891 (.a(n_3619), .y(add_88_69_n_1741));
nand2 add_88_69_g1892 (.a(n_1217), .b(n_3502), .y(add_88_69_n_1743));
nand2 add_88_69_g1893 (.a(n_1239), .b(n_1244), .y(add_88_69_n_1745));
nand2 add_88_69_g1894 (.a(n_968), .b(n_3611), .y(add_88_69_n_1746));
nand2 add_88_69_g1895 (.a(n_988), .b(n_3139), .y(add_88_69_n_1749));
nand2 add_88_69_g1896 (.a(n_3707), .b(n_3272), .y(add_88_69_n_1702));
nand2 add_88_69_g1897 (.a(n_1241), .b(n_1246), .y(add_88_69_n_1703));
nand2 add_88_69_g1898 (.a(n_3914), .b(n_3611), .y(add_88_69_n_1705));
nand2 add_88_69_g1900 (.a(n_3712), .b(n_2005), .y(add_88_69_n_1709));
nand2 add_88_69_g1901 (.a(n_2731), .b(n_3580), .y(add_88_69_n_1752));
nand2 add_88_69_g1902 (.a(n_986), .b(n_1240), .y(add_88_69_n_1755));
nor2 add_88_69_g1904 (.a(n_3707), .b(n_3272), .y(add_88_69_n_1714));
nor2 add_88_69_g1905 (.a(n_3914), .b(n_3611), .y(add_88_69_n_1716));
nand2 add_88_69_g1906 (.a(n_967), .b(n_3502), .y(add_88_69_n_1717));
nor2 add_88_69_g1907 (.a(n_1239), .b(n_1244), .y(add_88_69_n_1718));
nor2 add_88_69_g1908 (.a(n_3712), .b(n_2005), .y(add_88_69_n_1720));
nor2 add_88_69_g1909 (.a(n_985), .b(n_1239), .y(add_88_69_n_1722));
nand2 add_88_69_g1910 (.a(n_985), .b(n_1239), .y(add_88_69_n_1723));
nand2 add_88_69_g1913 (.a(n_3271), .b(n_1243), .y(add_88_69_n_1728));
nor2 add_88_69_g1914 (.a(n_1240), .b(n_1245), .y(add_88_69_n_1729));
nor2 add_88_69_g1915 (.a(n_3271), .b(n_1243), .y(add_88_69_n_1731));
nand2 add_88_69_g1917 (.a(n_2194), .b(n_3708), .y(add_88_69_n_1735));
nor2 add_88_69_g1918 (.a(n_981), .b(n_1235), .y(add_88_69_n_1737));
nor2 add_88_69_g1920 (.a(n_3607), .b(n_2033), .y(add_88_69_n_1739));
nor2 add_88_69_g1921 (.a(n_975), .b(n_4048), .y(add_88_69_n_1740));
xor2 add_88_21_g1052 (.a(n_3284), .b(add_88_21_n_1005), .y(n_736));
inv add_88_21_g1060 (.a(n_3894), .y(add_88_21_n_673));
nor2 add_88_21_g1066 (.a(n_2135), .b(n_3284), .y(add_88_21_n_681));
nand2 add_88_21_g1073 (.a(n_1313), .b(add_88_21_n_693), .y(add_88_21_n_688));
inv add_88_21_g1077 (.a(n_3284), .y(add_88_21_n_693));
xor2 add_88_21_g1095 (.a(add_88_21_n_726), .b(add_88_21_n_1012), .y(n_728));
nor2 add_88_21_g1097 (.a(add_88_21_n_726), .b(add_88_21_n_871), .y(add_88_21_n_713));
inv add_88_21_g1098 (.a(add_88_21_n_716), .y(add_88_21_n_715));
nor2 add_88_21_g1099 (.a(add_88_21_n_726), .b(add_88_21_n_1108), .y(add_88_21_n_716));
nand2 add_88_21_g1101 (.a(add_88_21_n_727), .b(add_88_21_n_923), .y(add_88_21_n_718));
nor2 add_88_21_g1102 (.a(add_88_21_n_845), .b(add_88_21_n_726), .y(add_88_21_n_720));
nor2 add_88_21_g1103 (.a(add_88_21_n_726), .b(add_88_21_n_907), .y(add_88_21_n_721));
inv add_88_21_g1108 (.a(add_88_21_n_726), .y(add_88_21_n_727));
nor2 add_88_21_g1109 (.a(add_88_21_n_795), .b(add_88_21_n_735), .y(add_88_21_n_726));
nor2 add_88_21_g1113 (.a(add_88_21_n_746), .b(add_88_21_n_1133), .y(add_88_21_n_731));
nor2 add_88_21_g1114 (.a(add_88_21_n_753), .b(n_3325), .y(add_88_21_n_733));
nand2 add_88_21_g1115 (.a(add_88_21_n_747), .b(add_88_21_n_929), .y(add_88_21_n_734));
nor2 add_88_21_g1116 (.a(add_88_21_n_919), .b(add_88_21_n_753), .y(add_88_21_n_735));
nand2 add_88_21_g1120 (.a(add_88_21_n_747), .b(add_88_21_n_843), .y(add_88_21_n_741));
nor2 add_88_21_g1121 (.a(add_88_21_n_746), .b(n_3891), .y(add_88_21_n_742));
nor2 add_88_21_g1122 (.a(add_88_21_n_746), .b(add_88_21_n_841), .y(add_88_21_n_743));
nand2 add_88_21_g1123 (.a(add_88_21_n_747), .b(add_88_21_n_869), .y(add_88_21_n_744));
xor2 add_88_21_g1124 (.a(add_88_21_n_997), .b(add_88_21_n_771), .y(n_724));
inv add_88_21_g1125 (.a(add_88_21_n_746), .y(add_88_21_n_747));
nor2 add_88_21_g1127 (.a(add_88_21_n_768), .b(add_88_21_n_1055), .y(add_88_21_n_749));
nand2 add_88_21_g1128 (.a(add_88_21_n_760), .b(add_88_21_n_874), .y(add_88_21_n_750));
nand2 add_88_21_g1129 (.a(add_88_21_n_762), .b(add_88_21_n_901), .y(add_88_21_n_751));
nor2 add_88_21_g1131 (.a(add_88_21_n_799), .b(add_88_21_n_769), .y(add_88_21_n_746));
nand2 add_88_21_g1134 (.a(add_88_21_n_771), .b(add_88_21_n_1062), .y(add_88_21_n_756));
nand2 add_88_21_g1135 (.a(add_88_21_n_783), .b(add_88_21_n_775), .y(add_88_21_n_758));
nand2 add_88_21_g1137 (.a(add_88_21_n_953), .b(add_88_21_n_771), .y(add_88_21_n_753));
nand2 add_88_21_g1138 (.a(add_88_21_n_778), .b(add_88_21_n_925), .y(add_88_21_n_760));
nand2 add_88_21_g1139 (.a(add_88_21_n_781), .b(add_88_21_n_927), .y(add_88_21_n_762));
nand2 add_88_21_g1140 (.a(add_88_21_n_797), .b(n_2853), .y(add_88_21_n_764));
nor2 add_88_21_g1142 (.a(add_88_21_n_779), .b(n_1591), .y(add_88_21_n_768));
nor2 add_88_21_g1143 (.a(add_88_21_n_779), .b(add_88_21_n_865), .y(add_88_21_n_769));
nor2 add_88_21_g1144 (.a(add_88_21_n_780), .b(add_88_21_n_1132), .y(add_88_21_n_772));
nor2 add_88_21_g1145 (.a(add_88_21_n_796), .b(add_88_21_n_895), .y(add_88_21_n_773));
nand2 add_88_21_g1146 (.a(add_88_21_n_797), .b(n_2854), .y(add_88_21_n_774));
nand2 add_88_21_g1147 (.a(add_88_21_n_778), .b(add_88_21_n_866), .y(add_88_21_n_775));
nand2 add_88_21_g1149 (.a(add_88_21_n_911), .b(add_88_21_n_1256), .y(add_88_21_n_771));
inv add_88_21_g1150 (.a(add_88_21_n_778), .y(add_88_21_n_779));
inv add_88_21_g1151 (.a(add_88_21_n_781), .y(add_88_21_n_780));
nor2 add_88_21_g1152 (.a(add_88_21_n_834), .b(add_88_21_n_1039), .y(add_88_21_n_783));
nor2 add_88_21_g1154 (.a(add_88_21_n_826), .b(add_88_21_n_1060), .y(add_88_21_n_787));
nand2 add_88_21_g1155 (.a(add_88_21_n_838), .b(add_88_21_n_1117), .y(add_88_21_n_788));
nor2 add_88_21_g1156 (.a(n_1316), .b(add_88_21_n_1133), .y(add_88_21_n_789));
nand2 add_88_21_g1157 (.a(n_2846), .b(add_88_21_n_929), .y(add_88_21_n_791));
nand2 add_88_21_g1158 (.a(add_88_21_n_813), .b(n_1598), .y(add_88_21_n_793));
nand2 add_88_21_g1160 (.a(add_88_21_n_903), .b(add_88_21_n_856), .y(add_88_21_n_795));
nand2 add_88_21_g1161 (.a(add_88_21_n_904), .b(add_88_21_n_847), .y(add_88_21_n_778));
nand2 add_88_21_g1162 (.a(add_88_21_n_833), .b(add_88_21_n_884), .y(add_88_21_n_781));
inv add_88_21_g1163 (.a(add_88_21_n_797), .y(add_88_21_n_796));
nand2 add_88_21_g1164 (.a(add_88_21_n_819), .b(add_88_21_n_909), .y(add_88_21_n_799));
nand2 add_88_21_g1165 (.a(add_88_21_n_848), .b(n_3423), .y(add_88_21_n_800));
nand2 add_88_21_g1166 (.a(add_88_21_n_839), .b(n_3326), .y(add_88_21_n_801));
xor2 add_88_21_g1167 (.a(add_88_21_n_1022), .b(add_88_21_n_876), .y(n_722));
nand2 add_88_21_g1168 (.a(n_2846), .b(add_88_21_n_869), .y(add_88_21_n_803));
nand2 add_88_21_g1169 (.a(add_88_21_n_859), .b(add_88_21_n_910), .y(add_88_21_n_805));
nand2 add_88_21_g1170 (.a(add_88_21_n_840), .b(n_1804), .y(add_88_21_n_806));
nor2 add_88_21_g1173 (.a(n_3891), .b(n_1316), .y(add_88_21_n_810));
nand2 add_88_21_g1174 (.a(add_88_21_n_815), .b(n_3170), .y(add_88_21_n_812));
nand2 add_88_21_g1175 (.a(add_88_21_n_905), .b(add_88_21_n_825), .y(add_88_21_n_797));
inv add_88_21_g1176 (.a(add_88_21_n_823), .y(add_88_21_n_813));
nand2 add_88_21_g1179 (.a(add_88_21_n_875), .b(add_88_21_n_916), .y(add_88_21_n_819));
nor2 add_88_21_g1180 (.a(add_88_21_n_882), .b(n_1591), .y(add_88_21_n_820));
nor2 add_88_21_g1181 (.a(add_88_21_n_872), .b(n_1597), .y(add_88_21_n_823));
nand2 add_88_21_g1182 (.a(add_88_21_n_917), .b(add_88_21_n_898), .y(add_88_21_n_825));
nor2 add_88_21_g1183 (.a(add_88_21_n_897), .b(n_2118), .y(add_88_21_n_826));
nand2 add_88_21_g1184 (.a(add_88_21_n_883), .b(add_88_21_n_925), .y(add_88_21_n_828));
nor2 add_88_21_g1185 (.a(add_88_21_n_871), .b(add_88_21_n_1132), .y(add_88_21_n_830));
nand2 add_88_21_g1186 (.a(add_88_21_n_878), .b(add_88_21_n_915), .y(add_88_21_n_833));
nor2 add_88_21_g1187 (.a(add_88_21_n_874), .b(n_3726), .y(add_88_21_n_834));
nand2 add_88_21_g1188 (.a(add_88_21_n_1103), .b(add_88_21_n_876), .y(add_88_21_n_815));
inv add_88_21_g1191 (.a(add_88_21_n_850), .y(add_88_21_n_838));
inv add_88_21_g1192 (.a(add_88_21_n_852), .y(add_88_21_n_839));
inv add_88_21_g1193 (.a(add_88_21_n_857), .y(add_88_21_n_840));
inv add_88_21_g1194 (.a(n_2136), .y(add_88_21_n_841));
inv add_88_21_g1195 (.a(n_1315), .y(add_88_21_n_843));
nand2 add_88_21_g1196 (.a(add_88_21_n_927), .b(add_88_21_n_870), .y(add_88_21_n_845));
nand2 add_88_21_g1197 (.a(add_88_21_n_921), .b(add_88_21_n_873), .y(add_88_21_n_847));
nand2 add_88_21_g1198 (.a(add_88_21_n_878), .b(add_88_21_n_1072), .y(add_88_21_n_848));
nor2 add_88_21_g1199 (.a(add_88_21_n_901), .b(add_88_21_n_1139), .y(add_88_21_n_850));
nor2 add_88_21_g1200 (.a(add_88_21_n_900), .b(n_3325), .y(add_88_21_n_852));
xor2 add_88_21_g1201 (.a(add_88_21_n_985), .b(n_3145), .y(n_721));
nand2 add_88_21_g1202 (.a(add_88_21_n_920), .b(add_88_21_n_899), .y(add_88_21_n_856));
nor2 add_88_21_g1203 (.a(add_88_21_n_868), .b(n_1805), .y(add_88_21_n_857));
nand2 add_88_21_g1204 (.a(add_88_21_n_902), .b(add_88_21_n_918), .y(add_88_21_n_859));
nand2 add_88_21_g1205 (.a(add_88_21_n_866), .b(add_88_21_n_883), .y(add_88_21_n_860));
inv add_88_21_g1209 (.a(add_88_21_n_871), .y(add_88_21_n_870));
inv add_88_21_g1210 (.a(add_88_21_n_872), .y(add_88_21_n_873));
inv add_88_21_g1211 (.a(add_88_21_n_874), .y(add_88_21_n_875));
inv add_88_21_g1212 (.a(add_88_21_n_878), .y(add_88_21_n_877));
inv add_88_21_g1214 (.a(add_88_21_n_882), .y(add_88_21_n_883));
nor2 add_88_21_g1215 (.a(add_88_21_n_939), .b(add_88_21_n_1024), .y(add_88_21_n_884));
nand2 add_88_21_g1216 (.a(add_88_21_n_916), .b(add_88_21_n_925), .y(add_88_21_n_865));
nor2 add_88_21_g1217 (.a(add_88_21_n_926), .b(n_3726), .y(add_88_21_n_866));
nand2 add_88_21_g1218 (.a(add_88_21_n_918), .b(add_88_21_n_927), .y(add_88_21_n_887));
nor2 add_88_21_g1219 (.a(add_88_21_n_944), .b(add_88_21_n_1033), .y(add_88_21_n_868));
nor2 add_88_21_g1220 (.a(n_2118), .b(add_88_21_n_930), .y(add_88_21_n_869));
nand2 add_88_21_g1221 (.a(add_88_21_n_915), .b(add_88_21_n_923), .y(add_88_21_n_871));
nor2 add_88_21_g1222 (.a(add_88_21_n_937), .b(add_88_21_n_1032), .y(add_88_21_n_872));
nor2 add_88_21_g1223 (.a(add_88_21_n_941), .b(add_88_21_n_1030), .y(add_88_21_n_874));
nand2 add_88_21_g1224 (.a(add_88_21_n_913), .b(n_3163), .y(add_88_21_n_876));
nand2 add_88_21_g1225 (.a(add_88_21_n_914), .b(n_3279), .y(add_88_21_n_878));
nand2 add_88_21_g1227 (.a(add_88_21_n_921), .b(add_88_21_n_924), .y(add_88_21_n_882));
inv add_88_21_g1228 (.a(add_88_21_n_897), .y(add_88_21_n_898));
inv add_88_21_g1229 (.a(add_88_21_n_900), .y(add_88_21_n_899));
inv add_88_21_g1230 (.a(add_88_21_n_901), .y(add_88_21_n_902));
nor2 add_88_21_g1231 (.a(add_88_21_n_947), .b(add_88_21_n_1037), .y(add_88_21_n_903));
nor2 add_88_21_g1232 (.a(add_88_21_n_949), .b(add_88_21_n_1028), .y(add_88_21_n_904));
nor2 add_88_21_g1233 (.a(add_88_21_n_933), .b(add_88_21_n_1026), .y(add_88_21_n_905));
nand2 add_88_21_g1234 (.a(add_88_21_n_1134), .b(add_88_21_n_924), .y(add_88_21_n_906));
nand2 add_88_21_g1235 (.a(add_88_21_n_923), .b(add_88_21_n_1072), .y(add_88_21_n_907));
nor2 add_88_21_g1236 (.a(add_88_21_n_957), .b(add_88_21_n_1095), .y(add_88_21_n_909));
nor2 add_88_21_g1237 (.a(add_88_21_n_931), .b(add_88_21_n_1097), .y(add_88_21_n_910));
nor2 add_88_21_g1238 (.a(add_88_21_n_955), .b(add_88_21_n_1093), .y(add_88_21_n_911));
nand2 add_88_21_g1239 (.a(n_2853), .b(n_1806), .y(add_88_21_n_895));
nor2 add_88_21_g1240 (.a(add_88_21_n_928), .b(add_88_21_n_1139), .y(add_88_21_n_896));
nor2 add_88_21_g1241 (.a(add_88_21_n_946), .b(n_1732), .y(add_88_21_n_897));
nor2 add_88_21_g1242 (.a(add_88_21_n_951), .b(add_88_21_n_1099), .y(add_88_21_n_900));
nor2 add_88_21_g1243 (.a(add_88_21_n_934), .b(add_88_21_n_1023), .y(add_88_21_n_901));
inv add_88_21_g1244 (.a(add_88_21_n_935), .y(add_88_21_n_913));
inv add_88_21_g1245 (.a(add_88_21_n_942), .y(add_88_21_n_914));
inv add_88_21_g1246 (.a(add_88_21_n_920), .y(add_88_21_n_919));
inv add_88_21_g1247 (.a(add_88_21_n_925), .y(add_88_21_n_926));
inv add_88_21_g1248 (.a(add_88_21_n_927), .y(add_88_21_n_928));
inv add_88_21_g1249 (.a(add_88_21_n_929), .y(add_88_21_n_930));
nor2 add_88_21_g1250 (.a(add_88_21_n_1112), .b(add_88_21_n_1117), .y(add_88_21_n_931));
nor2 add_88_21_g1251 (.a(n_1742), .b(n_2201), .y(add_88_21_n_933));
nor2 add_88_21_g1252 (.a(n_3404), .b(add_88_21_n_1053), .y(add_88_21_n_934));
nor2 add_88_21_g1253 (.a(n_3162), .b(n_3145), .y(add_88_21_n_935));
nor2 add_88_21_g1254 (.a(n_1624), .b(add_88_21_n_1126), .y(add_88_21_n_937));
nor2 add_88_21_g1255 (.a(n_3423), .b(n_3367), .y(add_88_21_n_939));
nor2 add_88_21_g1256 (.a(n_1590), .b(n_3299), .y(add_88_21_n_941));
nor2 add_88_21_g1257 (.a(n_3278), .b(add_88_21_n_1113), .y(add_88_21_n_942));
nor2 add_88_21_g1258 (.a(n_1782), .b(n_2125), .y(add_88_21_n_944));
nor2 add_88_21_g1259 (.a(n_1712), .b(add_88_21_n_1119), .y(add_88_21_n_946));
nor2 add_88_21_g1260 (.a(n_3336), .b(n_3326), .y(add_88_21_n_947));
nor2 add_88_21_g1261 (.a(n_1598), .b(n_3292), .y(add_88_21_n_949));
nor2 add_88_21_g1262 (.a(n_3191), .b(add_88_21_n_1042), .y(add_88_21_n_951));
nor2 add_88_21_g1263 (.a(n_3191), .b(add_88_21_n_1063), .y(add_88_21_n_953));
nor2 add_88_21_g1264 (.a(n_3184), .b(n_3170), .y(add_88_21_n_955));
nor2 add_88_21_g1265 (.a(n_1584), .b(n_3637), .y(add_88_21_n_957));
nor2 add_88_21_g1266 (.a(n_3367), .b(n_3424), .y(add_88_21_n_915));
nor2 add_88_21_g1267 (.a(n_3637), .b(n_3726), .y(add_88_21_n_916));
nor2 add_88_21_g1270 (.a(n_2201), .b(n_2118), .y(add_88_21_n_917));
nor2 add_88_21_g1271 (.a(add_88_21_n_1112), .b(add_88_21_n_1139), .y(add_88_21_n_918));
nor2 add_88_21_g1272 (.a(n_3336), .b(n_3325), .y(add_88_21_n_920));
nor2 add_88_21_g1273 (.a(n_3292), .b(n_1597), .y(add_88_21_n_921));
nor2 add_88_21_g1275 (.a(n_3278), .b(add_88_21_n_1108), .y(add_88_21_n_923));
nor2 add_88_21_g1276 (.a(n_1624), .b(add_88_21_n_1123), .y(add_88_21_n_924));
nor2 add_88_21_g1277 (.a(n_3299), .b(n_1591), .y(add_88_21_n_925));
nor2 add_88_21_g1278 (.a(n_3404), .b(add_88_21_n_1132), .y(add_88_21_n_927));
nor2 add_88_21_g1279 (.a(n_1712), .b(add_88_21_n_1133), .y(add_88_21_n_929));
nand2 add_88_21_g1281 (.a(add_88_21_n_1117), .b(add_88_21_n_1138), .y(add_88_21_n_979));
nand2 add_88_21_g1282 (.a(n_1584), .b(add_88_21_n_1140), .y(add_88_21_n_980));
nor2 add_88_21_g1283 (.a(add_88_21_n_1093), .b(n_3184), .y(add_88_21_n_982));
nand2 add_88_21_g1284 (.a(n_3163), .b(add_88_21_n_1035), .y(add_88_21_n_985));
nor2 add_88_21_g1285 (.a(add_88_21_n_1099), .b(n_3191), .y(add_88_21_n_987));
nor2 add_88_21_g1286 (.a(add_88_21_n_1030), .b(n_3299), .y(add_88_21_n_989));
nand2 add_88_21_g1287 (.a(n_1393), .b(add_88_21_n_1064), .y(add_88_21_n_991));
nor2 add_88_21_g1288 (.a(add_88_21_n_1101), .b(n_3278), .y(add_88_21_n_992));
nand2 add_88_21_g1290 (.a(n_1544), .b(add_88_21_n_1050), .y(add_88_21_n_996));
nor2 add_88_21_g1291 (.a(add_88_21_n_1043), .b(add_88_21_n_1063), .y(add_88_21_n_997));
nand2 add_88_21_g1292 (.a(add_88_21_n_1098), .b(add_88_21_n_1111), .y(add_88_21_n_999));
nor2 add_88_21_g1293 (.a(add_88_21_n_1023), .b(n_3404), .y(add_88_21_n_1000));
nor2 add_88_21_g1294 (.a(add_88_21_n_1129), .b(n_1597), .y(add_88_21_n_1002));
nand2 add_88_21_g1295 (.a(n_1590), .b(add_88_21_n_1142), .y(add_88_21_n_1003));
nand2 add_88_21_g1296 (.a(add_88_21_n_1126), .b(add_88_21_n_1122), .y(add_88_21_n_1005));
nor2 add_88_21_g1297 (.a(add_88_21_n_1032), .b(n_1624), .y(add_88_21_n_1006));
nor2 add_88_21_g1298 (.a(add_88_21_n_1127), .b(n_3424), .y(add_88_21_n_1008));
nand2 add_88_21_g1299 (.a(add_88_21_n_1053), .b(add_88_21_n_1131), .y(add_88_21_n_1010));
nand2 add_88_21_g1300 (.a(add_88_21_n_1113), .b(add_88_21_n_1107), .y(add_88_21_n_1012));
nand2 add_88_21_g1301 (.a(n_3207), .b(add_88_21_n_1105), .y(add_88_21_n_1013));
nor2 add_88_21_g1302 (.a(add_88_21_n_1049), .b(n_3325), .y(add_88_21_n_1014));
nand2 add_88_21_g1303 (.a(n_3368), .b(add_88_21_n_1067), .y(add_88_21_n_1015));
nor2 add_88_21_g1308 (.a(add_88_21_n_1118), .b(add_88_21_n_1133), .y(add_88_21_n_1020));
nor2 add_88_21_g1309 (.a(add_88_21_n_1121), .b(n_3169), .y(add_88_21_n_1022));
inv add_88_21_g1310 (.a(n_3405), .y(add_88_21_n_1023));
inv add_88_21_g1311 (.a(n_3368), .y(add_88_21_n_1024));
inv add_88_21_g1312 (.a(n_1762), .y(add_88_21_n_1026));
inv add_88_21_g1313 (.a(n_1544), .y(add_88_21_n_1028));
inv add_88_21_g1314 (.a(n_1487), .y(add_88_21_n_1030));
inv add_88_21_g1316 (.a(n_1625), .y(add_88_21_n_1032));
inv add_88_21_g1317 (.a(n_1674), .y(add_88_21_n_1033));
inv add_88_21_g1318 (.a(n_3162), .y(add_88_21_n_1035));
inv add_88_21_g1319 (.a(n_3207), .y(add_88_21_n_1037));
inv add_88_21_g1320 (.a(n_1584), .y(add_88_21_n_1039));
inv add_88_21_g1321 (.a(add_88_21_n_1042), .y(add_88_21_n_1043));
inv add_88_21_g1323 (.a(n_3326), .y(add_88_21_n_1049));
inv add_88_21_g1324 (.a(n_3292), .y(add_88_21_n_1050));
inv add_88_21_g1326 (.a(n_1590), .y(add_88_21_n_1055));
inv add_88_21_g1329 (.a(add_88_21_n_1063), .y(add_88_21_n_1062));
inv add_88_21_g1330 (.a(n_3637), .y(add_88_21_n_1064));
inv add_88_21_g1331 (.a(n_3367), .y(add_88_21_n_1067));
inv add_88_21_g1333 (.a(n_3424), .y(add_88_21_n_1072));
nand2 add_88_21_g1346 (.a(n_764), .b(v1_4_), .y(add_88_21_n_1042));
nand2 add_88_21_g1352 (.a(n_788), .b(v1_12_), .y(add_88_21_n_1053));
nor2 add_88_21_g1358 (.a(n_764), .b(v1_4_), .y(add_88_21_n_1063));
inv add_88_21_g1364 (.a(n_3185), .y(add_88_21_n_1093));
inv add_88_21_g1365 (.a(n_1393), .y(add_88_21_n_1095));
inv add_88_21_g1366 (.a(add_88_21_n_1098), .y(add_88_21_n_1097));
inv add_88_21_g1367 (.a(n_3192), .y(add_88_21_n_1099));
inv add_88_21_g1368 (.a(n_3279), .y(add_88_21_n_1101));
inv add_88_21_g1369 (.a(n_3169), .y(add_88_21_n_1103));
inv add_88_21_g1370 (.a(n_3336), .y(add_88_21_n_1105));
inv add_88_21_g1371 (.a(add_88_21_n_1108), .y(add_88_21_n_1107));
inv add_88_21_g1373 (.a(add_88_21_n_1112), .y(add_88_21_n_1111));
inv add_88_21_g1375 (.a(add_88_21_n_1119), .y(add_88_21_n_1118));
inv add_88_21_g1376 (.a(n_3170), .y(add_88_21_n_1121));
inv add_88_21_g1377 (.a(add_88_21_n_1123), .y(add_88_21_n_1122));
inv add_88_21_g1379 (.a(n_3423), .y(add_88_21_n_1127));
inv add_88_21_g1380 (.a(n_1598), .y(add_88_21_n_1129));
inv add_88_21_g1381 (.a(add_88_21_n_1132), .y(add_88_21_n_1131));
inv add_88_21_g1382 (.a(n_1597), .y(add_88_21_n_1134));
inv add_88_21_g1384 (.a(add_88_21_n_1139), .y(add_88_21_n_1138));
inv add_88_21_g1385 (.a(n_3726), .y(add_88_21_n_1140));
inv add_88_21_g1386 (.a(n_1591), .y(add_88_21_n_1142));
nand2 add_88_21_g1390 (.a(n_797), .b(v1_15_), .y(add_88_21_n_1098));
nor2 add_88_21_g1396 (.a(n_776), .b(v1_8_), .y(add_88_21_n_1108));
nor2 add_88_21_g1398 (.a(n_797), .b(v1_15_), .y(add_88_21_n_1112));
nand2 add_88_21_g1399 (.a(n_776), .b(v1_8_), .y(add_88_21_n_1113));
nand2 add_88_21_g1402 (.a(n_794), .b(v1_14_), .y(add_88_21_n_1117));
nand2 add_88_21_g1403 (.a(n_2121), .b(v1_24_), .y(add_88_21_n_1119));
nor2 add_88_21_g1405 (.a(n_2197), .b(v1_16_), .y(add_88_21_n_1123));
nand2 add_88_21_g1407 (.a(n_2197), .b(v1_16_), .y(add_88_21_n_1126));
nor2 add_88_21_g1410 (.a(n_788), .b(v1_12_), .y(add_88_21_n_1132));
nor2 add_88_21_g1411 (.a(n_2121), .b(v1_24_), .y(add_88_21_n_1133));
nor2 add_88_21_g1414 (.a(n_794), .b(v1_14_), .y(add_88_21_n_1139));
inv add_88_21_g3 (.a(add_88_21_n_1255), .y(add_88_21_n_1256));
nor2 add_88_21_g2 (.a(n_3184), .b(add_88_21_n_815), .y(add_88_21_n_1255));
xor2 add_76_21_g1144 (.a(add_76_21_n_805), .b(add_76_21_n_1163), .y(n_1224));
xor2 add_76_21_g1146 (.a(add_76_21_n_799), .b(add_76_21_n_1160), .y(n_1216));
xor2 add_76_21_g1147 (.a(n_3733), .b(add_76_21_n_1161), .y(n_1217));
nand2 add_76_21_g1164 (.a(add_76_21_n_851), .b(n_3438), .y(add_76_21_n_799));
nand2 add_76_21_g1165 (.a(n_2833), .b(n_3941), .y(add_76_21_n_800));
nor2 add_76_21_g1169 (.a(add_76_21_n_824), .b(add_76_21_n_929), .y(add_76_21_n_804));
nor2 add_76_21_g1170 (.a(add_76_21_n_819), .b(add_76_21_n_888), .y(add_76_21_n_805));
nor2 add_76_21_g1175 (.a(n_3710), .b(add_76_21_n_919), .y(add_76_21_n_811));
nor2 add_76_21_g1178 (.a(n_3710), .b(add_76_21_n_926), .y(add_76_21_n_815));
nor2 add_76_21_g1180 (.a(n_3710), .b(add_76_21_n_961), .y(add_76_21_n_817));
nor2 add_76_21_g1181 (.a(n_3710), .b(add_76_21_n_1011), .y(add_76_21_n_818));
nor2 add_76_21_g1182 (.a(n_3710), .b(add_76_21_n_995), .y(add_76_21_n_819));
nor2 add_76_21_g1183 (.a(n_3710), .b(add_76_21_n_938), .y(add_76_21_n_820));
nor2 add_76_21_g1187 (.a(n_3710), .b(add_76_21_n_1044), .y(add_76_21_n_824));
xor2 add_76_21_g1191 (.a(add_76_21_n_835), .b(add_76_21_n_1137), .y(n_1235));
nor2 add_76_21_g1198 (.a(n_3662), .b(add_76_21_n_858), .y(add_76_21_n_835));
nand2 add_76_21_g1200 (.a(add_76_21_n_846), .b(n_2018), .y(add_76_21_n_837));
xor2 add_76_21_g1203 (.a(add_76_21_n_872), .b(add_76_21_n_1148), .y(n_1241));
xor2 add_76_21_g1204 (.a(add_76_21_n_878), .b(add_76_21_n_1127), .y(n_1240));
xor2 add_76_21_g1205 (.a(n_2946), .b(add_76_21_n_1130), .y(n_1239));
inv add_76_21_g1209 (.a(add_76_21_n_854), .y(add_76_21_n_846));
nor2 add_76_21_g1214 (.a(add_76_21_n_886), .b(add_76_21_n_875), .y(add_76_21_n_851));
nor2 add_76_21_g1216 (.a(n_2946), .b(n_4092), .y(add_76_21_n_854));
nor2 add_76_21_g1219 (.a(n_2946), .b(n_3700), .y(add_76_21_n_858));
nor2 add_76_21_g1220 (.a(add_76_21_n_988), .b(n_2946), .y(add_76_21_n_859));
nor2 add_76_21_g1222 (.a(add_76_21_n_992), .b(n_2946), .y(add_76_21_n_861));
nor2 add_76_21_g1224 (.a(n_2946), .b(n_2966), .y(add_76_21_n_863));
nand2 add_76_21_g1230 (.a(add_76_21_n_884), .b(add_76_21_n_1034), .y(add_76_21_n_872));
nor2 add_76_21_g1234 (.a(n_3941), .b(add_76_21_n_977), .y(add_76_21_n_875));
xor2 add_76_21_g1236 (.a(add_76_21_n_906), .b(add_76_21_n_1119), .y(n_1243));
nand2 add_76_21_g1237 (.a(add_76_21_n_935), .b(add_76_21_n_894), .y(add_76_21_n_878));
nor2 add_76_21_g1239 (.a(add_76_21_n_1020), .b(add_76_21_n_907), .y(add_76_21_n_881));
nand2 add_76_21_g1240 (.a(add_76_21_n_896), .b(add_76_21_n_1009), .y(add_76_21_n_882));
nand2 add_76_21_g1242 (.a(add_76_21_n_906), .b(add_76_21_n_1065), .y(add_76_21_n_884));
nand2 add_76_21_g1243 (.a(add_76_21_n_908), .b(add_76_21_n_936), .y(add_76_21_n_886));
nand2 add_76_21_g1246 (.a(add_76_21_n_918), .b(add_76_21_n_912), .y(add_76_21_n_888));
nand2 add_76_21_g1247 (.a(add_76_21_n_906), .b(add_76_21_n_1240), .y(add_76_21_n_889));
nand2 add_76_21_g1248 (.a(add_76_21_n_900), .b(add_76_21_n_1005), .y(add_76_21_n_890));
nor2 add_76_21_g1249 (.a(add_76_21_n_911), .b(n_1952), .y(add_76_21_n_891));
nand2 add_76_21_g1251 (.a(add_76_21_n_913), .b(add_76_21_n_925), .y(add_76_21_n_893));
nand2 add_76_21_g1252 (.a(add_76_21_n_1045), .b(add_76_21_n_906), .y(add_76_21_n_894));
xor2 add_76_21_g1253 (.a(add_76_21_n_1150), .b(add_76_21_n_947), .y(n_1244));
nand2 add_76_21_g1254 (.a(add_76_21_n_914), .b(add_76_21_n_1070), .y(add_76_21_n_896));
nand2 add_76_21_g1256 (.a(n_1948), .b(add_76_21_n_1063), .y(add_76_21_n_900));
nor2 add_76_21_g1257 (.a(add_76_21_n_915), .b(n_1551), .y(add_76_21_n_902));
nor2 add_76_21_g1259 (.a(n_3663), .b(n_2340), .y(add_76_21_n_905));
inv add_76_21_g1260 (.a(add_76_21_n_906), .y(add_76_21_n_907));
nand2 add_76_21_g1261 (.a(n_1948), .b(add_76_21_n_1032), .y(add_76_21_n_908));
nor2 add_76_21_g1263 (.a(add_76_21_n_932), .b(n_3010), .y(add_76_21_n_911));
nand2 add_76_21_g1264 (.a(add_76_21_n_914), .b(add_76_21_n_1006), .y(add_76_21_n_912));
nand2 add_76_21_g1265 (.a(n_3662), .b(add_76_21_n_1031), .y(add_76_21_n_913));
nand2 add_76_21_g1266 (.a(add_76_21_n_1043), .b(add_76_21_n_1395), .y(add_76_21_n_906));
inv add_76_21_g1267 (.a(add_76_21_n_914), .y(add_76_21_n_915));
nor2 add_76_21_g1269 (.a(add_76_21_n_971), .b(add_76_21_n_1183), .y(add_76_21_n_918));
nand2 add_76_21_g1270 (.a(add_76_21_n_948), .b(add_76_21_n_949), .y(add_76_21_n_919));
nor2 add_76_21_g1271 (.a(add_76_21_n_964), .b(add_76_21_n_1185), .y(add_76_21_n_922));
nor2 add_76_21_g1273 (.a(add_76_21_n_990), .b(add_76_21_n_1195), .y(add_76_21_n_925));
nand2 add_76_21_g1274 (.a(add_76_21_n_949), .b(add_76_21_n_1072), .y(add_76_21_n_926));
nor2 add_76_21_g1275 (.a(add_76_21_n_959), .b(add_76_21_n_1017), .y(add_76_21_n_928));
nand2 add_76_21_g1276 (.a(add_76_21_n_975), .b(n_4499), .y(add_76_21_n_929));
nand2 add_76_21_g1277 (.a(add_76_21_n_984), .b(add_76_21_n_1041), .y(add_76_21_n_930));
nand2 add_76_21_g1278 (.a(add_76_21_n_1042), .b(add_76_21_n_985), .y(add_76_21_n_914));
nor2 add_76_21_g1283 (.a(add_76_21_n_968), .b(add_76_21_n_1263), .y(add_76_21_n_935));
nor2 add_76_21_g1284 (.a(add_76_21_n_966), .b(add_76_21_n_1172), .y(add_76_21_n_936));
xor2 add_76_21_g1285 (.a(add_76_21_n_1124), .b(add_76_21_n_1033), .y(n_1245));
nand2 add_76_21_g1286 (.a(add_76_21_n_949), .b(add_76_21_n_1004), .y(add_76_21_n_938));
nand2 add_76_21_g1287 (.a(n_4398), .b(n_1428), .y(add_76_21_n_940));
nor2 add_76_21_g1289 (.a(add_76_21_n_978), .b(add_76_21_n_950), .y(add_76_21_n_942));
nand2 add_76_21_g1291 (.a(add_76_21_n_980), .b(n_4356), .y(add_76_21_n_947));
inv add_76_21_g1293 (.a(add_76_21_n_949), .y(add_76_21_n_950));
nor2 add_76_21_g1294 (.a(n_3700), .b(n_2340), .y(add_76_21_n_951));
nor2 add_76_21_g1296 (.a(add_76_21_n_1002), .b(n_3700), .y(add_76_21_n_957));
nor2 add_76_21_g1297 (.a(add_76_21_n_1040), .b(add_76_21_n_1059), .y(add_76_21_n_959));
nand2 add_76_21_g1298 (.a(add_76_21_n_1012), .b(add_76_21_n_1070), .y(add_76_21_n_961));
nand2 add_76_21_g1299 (.a(add_76_21_n_1010), .b(add_76_21_n_1058), .y(add_76_21_n_963));
nor2 add_76_21_g1300 (.a(add_76_21_n_1038), .b(n_1662), .y(add_76_21_n_964));
nor2 add_76_21_g1301 (.a(add_76_21_n_1005), .b(add_76_21_n_1194), .y(add_76_21_n_966));
nor2 add_76_21_g1302 (.a(add_76_21_n_1034), .b(n_1512), .y(add_76_21_n_968));
nor2 add_76_21_g1304 (.a(add_76_21_n_1009), .b(n_1637), .y(add_76_21_n_971));
nor2 add_76_21_g1305 (.a(add_76_21_n_1015), .b(n_3010), .y(add_76_21_n_948));
nor2 add_76_21_g1306 (.a(add_76_21_n_1003), .b(add_76_21_n_1011), .y(add_76_21_n_949));
inv add_76_21_g1307 (.a(add_76_21_n_982), .y(add_76_21_n_975));
nand2 add_76_21_g1310 (.a(add_76_21_n_1039), .b(add_76_21_n_1056), .y(add_76_21_n_981));
nor2 add_76_21_g1311 (.a(n_4289), .b(n_3881), .y(add_76_21_n_982));
nand2 add_76_21_g1312 (.a(add_76_21_n_1035), .b(add_76_21_n_1057), .y(add_76_21_n_984));
nand2 add_76_21_g1313 (.a(n_4290), .b(add_76_21_n_1055), .y(add_76_21_n_985));
nand2 add_76_21_g1315 (.a(add_76_21_n_1014), .b(add_76_21_n_1068), .y(add_76_21_n_988));
nor2 add_76_21_g1316 (.a(add_76_21_n_1040), .b(n_2288), .y(add_76_21_n_990));
xor2 add_76_21_g1317 (.a(add_76_21_n_1117), .b(add_76_21_n_1192), .y(n_1246));
nand2 add_76_21_g1318 (.a(add_76_21_n_1031), .b(add_76_21_n_1014), .y(add_76_21_n_992));
nand2 add_76_21_g1319 (.a(add_76_21_n_1006), .b(add_76_21_n_1012), .y(add_76_21_n_995));
nand2 add_76_21_g1320 (.a(add_76_21_n_1032), .b(add_76_21_n_1016), .y(add_76_21_n_977));
nand2 add_76_21_g1321 (.a(add_76_21_n_1016), .b(add_76_21_n_1063), .y(add_76_21_n_978));
nand2 add_76_21_g1322 (.a(add_76_21_n_1033), .b(add_76_21_n_1231), .y(add_76_21_n_980));
inv add_76_21_g1324 (.a(add_76_21_n_1009), .y(add_76_21_n_1010));
inv add_76_21_g1325 (.a(add_76_21_n_1011), .y(add_76_21_n_1012));
inv add_76_21_g1326 (.a(n_3700), .y(add_76_21_n_1014));
inv add_76_21_g1327 (.a(add_76_21_n_1015), .y(add_76_21_n_1016));
nand2 add_76_21_g1328 (.a(add_76_21_n_1078), .b(n_1400), .y(add_76_21_n_1017));
nor2 add_76_21_g1329 (.a(add_76_21_n_1075), .b(add_76_21_n_1176), .y(add_76_21_n_1018));
nor2 add_76_21_g1330 (.a(add_76_21_n_1083), .b(add_76_21_n_1178), .y(add_76_21_n_1019));
nand2 add_76_21_g1331 (.a(add_76_21_n_1057), .b(add_76_21_n_1065), .y(add_76_21_n_1020));
nand2 add_76_21_g1332 (.a(add_76_21_n_1060), .b(add_76_21_n_1068), .y(add_76_21_n_1002));
nand2 add_76_21_g1333 (.a(add_76_21_n_1058), .b(add_76_21_n_1070), .y(add_76_21_n_1003));
nor2 add_76_21_g1334 (.a(add_76_21_n_1071), .b(n_1662), .y(add_76_21_n_1004));
nor2 add_76_21_g1335 (.a(add_76_21_n_1088), .b(add_76_21_n_1174), .y(add_76_21_n_1005));
nor2 add_76_21_g1336 (.a(add_76_21_n_1069), .b(n_1637), .y(add_76_21_n_1006));
nor2 add_76_21_g1338 (.a(add_76_21_n_1093), .b(add_76_21_n_1238), .y(add_76_21_n_1009));
nand2 add_76_21_g1339 (.a(add_76_21_n_1055), .b(n_1885), .y(add_76_21_n_1011));
nand2 add_76_21_g1341 (.a(add_76_21_n_1056), .b(add_76_21_n_1072), .y(add_76_21_n_1015));
inv add_76_21_g1342 (.a(add_76_21_n_1034), .y(add_76_21_n_1035));
inv add_76_21_g1344 (.a(add_76_21_n_1038), .y(add_76_21_n_1039));
nor2 add_76_21_g1345 (.a(add_76_21_n_1085), .b(add_76_21_n_1173), .y(add_76_21_n_1041));
nor2 add_76_21_g1346 (.a(n_3861), .b(add_76_21_n_1167), .y(add_76_21_n_1042));
nor2 add_76_21_g1347 (.a(add_76_21_n_1080), .b(add_76_21_n_1237), .y(add_76_21_n_1043));
nand2 add_76_21_g1348 (.a(n_1885), .b(add_76_21_n_1209), .y(add_76_21_n_1044));
nor2 add_76_21_g1349 (.a(add_76_21_n_1064), .b(n_1512), .y(add_76_21_n_1045));
nor2 add_76_21_g1350 (.a(add_76_21_n_1074), .b(add_76_21_n_1165), .y(add_76_21_n_1047));
nor2 add_76_21_g1352 (.a(add_76_21_n_1067), .b(n_2288), .y(add_76_21_n_1031));
nor2 add_76_21_g1353 (.a(add_76_21_n_1062), .b(add_76_21_n_1194), .y(add_76_21_n_1032));
nand2 add_76_21_g1354 (.a(add_76_21_n_1052), .b(n_3131), .y(add_76_21_n_1033));
nor2 add_76_21_g1355 (.a(n_2922), .b(add_76_21_n_1235), .y(add_76_21_n_1034));
nor2 add_76_21_g1357 (.a(add_76_21_n_1073), .b(n_1922), .y(add_76_21_n_1038));
nor2 add_76_21_g1358 (.a(add_76_21_n_1082), .b(add_76_21_n_1230), .y(add_76_21_n_1040));
inv add_76_21_g1359 (.a(add_76_21_n_1086), .y(add_76_21_n_1052));
inv add_76_21_g1361 (.a(add_76_21_n_1060), .y(add_76_21_n_1059));
inv add_76_21_g1362 (.a(add_76_21_n_1063), .y(add_76_21_n_1062));
inv add_76_21_g1363 (.a(add_76_21_n_1065), .y(add_76_21_n_1064));
inv add_76_21_g1364 (.a(add_76_21_n_1068), .y(add_76_21_n_1067));
inv add_76_21_g1365 (.a(add_76_21_n_1070), .y(add_76_21_n_1069));
inv add_76_21_g1366 (.a(add_76_21_n_1072), .y(add_76_21_n_1071));
nor2 add_76_21_g1367 (.a(n_1927), .b(n_2310), .y(add_76_21_n_1073));
nor2 add_76_21_g1368 (.a(n_1638), .b(n_1563), .y(add_76_21_n_1074));
nor2 add_76_21_g1369 (.a(n_1663), .b(n_3522), .y(add_76_21_n_1075));
nand2 add_76_21_g1371 (.a(add_76_21_n_1195), .b(add_76_21_n_1181), .y(add_76_21_n_1078));
nor2 add_76_21_g1372 (.a(n_3318), .b(n_4356), .y(add_76_21_n_1080));
nor2 add_76_21_g1373 (.a(n_1414), .b(n_2299), .y(add_76_21_n_1082));
nor2 add_76_21_g1374 (.a(n_1428), .b(n_3691), .y(add_76_21_n_1083));
nor2 add_76_21_g1375 (.a(n_1511), .b(n_2717), .y(add_76_21_n_1085));
nor2 add_76_21_g1376 (.a(n_3130), .b(add_76_21_n_1192), .y(add_76_21_n_1086));
nor2 add_76_21_g1377 (.a(n_3011), .b(n_2049), .y(add_76_21_n_1088));
nor2 add_76_21_g1380 (.a(n_1550), .b(n_1322), .y(add_76_21_n_1093));
nor2 add_76_21_g1384 (.a(n_2563), .b(n_3881), .y(add_76_21_n_1055));
nor2 add_76_21_g1385 (.a(n_3522), .b(n_1662), .y(add_76_21_n_1056));
nor2 add_76_21_g1386 (.a(n_2717), .b(n_1512), .y(add_76_21_n_1057));
nor2 add_76_21_g1388 (.a(n_1563), .b(n_1637), .y(add_76_21_n_1058));
nor2 add_76_21_g1389 (.a(n_2277), .b(n_2288), .y(add_76_21_n_1060));
nor2 add_76_21_g1391 (.a(n_2049), .b(n_3010), .y(add_76_21_n_1063));
nor2 add_76_21_g1392 (.a(n_2693), .b(n_2926), .y(add_76_21_n_1065));
nor2 add_76_21_g1394 (.a(n_2299), .b(n_2340), .y(add_76_21_n_1068));
nor2 add_76_21_g1395 (.a(n_1322), .b(n_1551), .y(add_76_21_n_1070));
nor2 add_76_21_g1396 (.a(n_2310), .b(n_1605), .y(add_76_21_n_1072));
nand2 add_76_21_g1399 (.a(n_3131), .b(add_76_21_n_1170), .y(add_76_21_n_1117));
nor2 add_76_21_g1400 (.a(n_2923), .b(n_2926), .y(add_76_21_n_1119));
nand2 add_76_21_g1401 (.a(n_1330), .b(add_76_21_n_1242), .y(add_76_21_n_1121));
nor2 add_76_21_g1402 (.a(n_1946), .b(n_1605), .y(add_76_21_n_1122));
nor2 add_76_21_g1403 (.a(add_76_21_n_1200), .b(n_4355), .y(add_76_21_n_1124));
nor2 add_76_21_g1405 (.a(add_76_21_n_1173), .b(n_2717), .y(add_76_21_n_1127));
nand2 add_76_21_g1407 (.a(n_2018), .b(add_76_21_n_1256), .y(add_76_21_n_1130));
nand2 add_76_21_g1409 (.a(n_1407), .b(add_76_21_n_1207), .y(add_76_21_n_1134));
nor2 add_76_21_g1410 (.a(add_76_21_n_1230), .b(n_2299), .y(add_76_21_n_1135));
nand2 add_76_21_g1411 (.a(n_1414), .b(add_76_21_n_1274), .y(add_76_21_n_1137));
nor2 add_76_21_g1413 (.a(add_76_21_n_1233), .b(n_3694), .y(add_76_21_n_1141));
nor2 add_76_21_g1415 (.a(add_76_21_n_1267), .b(n_3689), .y(add_76_21_n_1144));
nor2 add_76_21_g1417 (.a(add_76_21_n_1263), .b(n_1512), .y(add_76_21_n_1148));
nor2 add_76_21_g1418 (.a(add_76_21_n_1237), .b(n_3318), .y(add_76_21_n_1150));
nand2 add_76_21_g1420 (.a(n_3989), .b(add_76_21_n_1251), .y(add_76_21_n_1155));
nand2 add_76_21_g1421 (.a(n_4292), .b(add_76_21_n_1261), .y(add_76_21_n_1156));
nor2 add_76_21_g1423 (.a(add_76_21_n_1235), .b(n_2693), .y(add_76_21_n_1158));
xor2 add_76_21_g1424 (.a(n_941), .b(v0_31_), .y(add_76_21_n_1160));
nor2 add_76_21_g1425 (.a(add_76_21_n_1172), .b(add_76_21_n_1194), .y(add_76_21_n_1161));
nand2 add_76_21_g1426 (.a(n_1564), .b(add_76_21_n_1244), .y(add_76_21_n_1163));
inv add_76_21_g1427 (.a(n_1564), .y(add_76_21_n_1165));
inv add_76_21_g1428 (.a(n_1330), .y(add_76_21_n_1167));
inv add_76_21_g1430 (.a(n_3130), .y(add_76_21_n_1170));
inv add_76_21_g1431 (.a(add_76_21_n_1216), .y(add_76_21_n_1172));
inv add_76_21_g1432 (.a(n_1442), .y(add_76_21_n_1173));
inv add_76_21_g1433 (.a(n_3989), .y(add_76_21_n_1174));
inv add_76_21_g1434 (.a(n_3521), .y(add_76_21_n_1176));
inv add_76_21_g1435 (.a(n_1421), .y(add_76_21_n_1178));
inv add_76_21_g1436 (.a(n_2277), .y(add_76_21_n_1181));
inv add_76_21_g1437 (.a(n_1638), .y(add_76_21_n_1183));
inv add_76_21_g1438 (.a(n_1663), .y(add_76_21_n_1185));
inv add_76_21_g1441 (.a(n_1407), .y(add_76_21_n_1195));
inv add_76_21_g1443 (.a(n_4356), .y(add_76_21_n_1200));
inv add_76_21_g1445 (.a(n_1662), .y(add_76_21_n_1203));
inv add_76_21_g1447 (.a(n_2288), .y(add_76_21_n_1207));
nand2 add_76_21_g1454 (.a(n_938), .b(v0_30_), .y(add_76_21_n_1216));
nand2 add_76_21_g1466 (.a(n_848), .b(v0_0_), .y(add_76_21_n_1192));
nor2 add_76_21_g1468 (.a(n_938), .b(v0_30_), .y(add_76_21_n_1194));
inv add_76_21_g1479 (.a(n_1386), .y(add_76_21_n_1230));
inv add_76_21_g1480 (.a(n_4355), .y(add_76_21_n_1231));
inv add_76_21_g1481 (.a(n_2019), .y(add_76_21_n_1233));
inv add_76_21_g1482 (.a(n_1379), .y(add_76_21_n_1235));
inv add_76_21_g1484 (.a(n_3268), .y(add_76_21_n_1237));
inv add_76_21_g1485 (.a(n_1323), .y(add_76_21_n_1238));
inv add_76_21_g1486 (.a(n_2926), .y(add_76_21_n_1240));
inv add_76_21_g1487 (.a(n_2563), .y(add_76_21_n_1242));
inv add_76_21_g1488 (.a(n_1563), .y(add_76_21_n_1244));
inv add_76_21_g1490 (.a(n_1550), .y(add_76_21_n_1249));
inv add_76_21_g1491 (.a(n_2049), .y(add_76_21_n_1251));
inv add_76_21_g1492 (.a(n_3691), .y(add_76_21_n_1254));
inv add_76_21_g1493 (.a(n_4092), .y(add_76_21_n_1256));
inv add_76_21_g1495 (.a(n_1985), .y(add_76_21_n_1261));
inv add_76_21_g1496 (.a(n_1511), .y(add_76_21_n_1263));
inv add_76_21_g1497 (.a(n_1428), .y(add_76_21_n_1267));
inv add_76_21_g1499 (.a(n_1637), .y(add_76_21_n_1272));
inv add_76_21_g1500 (.a(n_2340), .y(add_76_21_n_1274));
inv add_76_21_g1501 (.a(n_1551), .y(add_76_21_n_1277));
inv add_76_21_g3 (.a(add_76_21_n_1394), .y(add_76_21_n_1395));
nor2 add_76_21_g2 (.a(n_3318), .b(add_76_21_n_980), .y(add_76_21_n_1394));
xor2 add_76_82_g1119 (.a(add_76_82_n_815), .b(add_76_82_n_1153), .y(n_939));
xor2 add_76_82_g1120 (.a(add_76_82_n_820), .b(add_76_82_n_1191), .y(n_942));
nand2 add_76_82_g1130 (.a(add_76_82_n_849), .b(add_76_82_n_854), .y(add_76_82_n_815));
nand2 add_76_82_g1135 (.a(add_76_82_n_842), .b(add_76_82_n_858), .y(add_76_82_n_820));
nor2 add_76_82_g1153 (.a(add_76_82_n_853), .b(add_76_82_n_949), .y(add_76_82_n_839));
nor2 add_76_82_g1154 (.a(add_76_82_n_853), .b(add_76_82_n_941), .y(add_76_82_n_840));
nand2 add_76_82_g1155 (.a(n_3866), .b(add_76_82_n_969), .y(add_76_82_n_842));
nor2 add_76_82_g1159 (.a(add_76_82_n_853), .b(add_76_82_n_984), .y(add_76_82_n_846));
nor2 add_76_82_g1160 (.a(add_76_82_n_853), .b(add_76_82_n_1040), .y(add_76_82_n_847));
nand2 add_76_82_g1161 (.a(n_3866), .b(add_76_82_n_1020), .y(add_76_82_n_848));
nand2 add_76_82_g1162 (.a(n_3866), .b(add_76_82_n_971), .y(add_76_82_n_849));
nand2 add_76_82_g1163 (.a(n_3866), .b(add_76_82_n_967), .y(add_76_82_n_850));
inv add_76_82_g1165 (.a(n_3866), .y(add_76_82_n_853));
nor2 add_76_82_g1166 (.a(add_76_82_n_895), .b(add_76_82_n_908), .y(add_76_82_n_854));
nand2 add_76_82_g1167 (.a(add_76_82_n_885), .b(add_76_82_n_909), .y(add_76_82_n_855));
nor2 add_76_82_g1168 (.a(add_76_82_n_888), .b(add_76_82_n_955), .y(add_76_82_n_856));
nor2 add_76_82_g1170 (.a(add_76_82_n_892), .b(add_76_82_n_905), .y(add_76_82_n_858));
nand2 add_76_82_g1176 (.a(add_76_82_n_879), .b(add_76_82_n_1063), .y(add_76_82_n_863));
nor2 add_76_82_g1177 (.a(add_76_82_n_893), .b(add_76_82_n_945), .y(add_76_82_n_864));
nand2 add_76_82_g1190 (.a(add_76_82_n_898), .b(add_76_82_n_1094), .y(add_76_82_n_879));
nand2 add_76_82_g1194 (.a(add_76_82_n_898), .b(add_76_82_n_976), .y(add_76_82_n_885));
nor2 add_76_82_g1196 (.a(n_2652), .b(add_76_82_n_1041), .y(add_76_82_n_888));
nor2 add_76_82_g1200 (.a(n_2652), .b(add_76_82_n_1004), .y(add_76_82_n_892));
nor2 add_76_82_g1201 (.a(n_2652), .b(add_76_82_n_1030), .y(add_76_82_n_893));
nor2 add_76_82_g1203 (.a(n_2652), .b(add_76_82_n_1005), .y(add_76_82_n_895));
inv add_76_82_g1204 (.a(n_2652), .y(add_76_82_n_898));
nor2 add_76_82_g1206 (.a(add_76_82_n_923), .b(add_76_82_n_1216), .y(add_76_82_n_901));
nor2 add_76_82_g1207 (.a(add_76_82_n_928), .b(add_76_82_n_1205), .y(add_76_82_n_902));
nand2 add_76_82_g1208 (.a(add_76_82_n_918), .b(add_76_82_n_1035), .y(add_76_82_n_903));
nand2 add_76_82_g1209 (.a(add_76_82_n_916), .b(add_76_82_n_1037), .y(add_76_82_n_904));
nand2 add_76_82_g1210 (.a(add_76_82_n_930), .b(add_76_82_n_961), .y(add_76_82_n_905));
nor2 add_76_82_g1211 (.a(add_76_82_n_922), .b(add_76_82_n_966), .y(add_76_82_n_896));
nand2 add_76_82_g1216 (.a(add_76_82_n_920), .b(add_76_82_n_1032), .y(add_76_82_n_908));
nor2 add_76_82_g1217 (.a(add_76_82_n_931), .b(add_76_82_n_1218), .y(add_76_82_n_909));
nor2 add_76_82_g1218 (.a(add_76_82_n_933), .b(add_76_82_n_940), .y(add_76_82_n_910));
nand2 add_76_82_g1219 (.a(add_76_82_n_934), .b(add_76_82_n_944), .y(add_76_82_n_911));
nor2 add_76_82_g1223 (.a(add_76_82_n_937), .b(add_76_82_n_1031), .y(add_76_82_n_915));
nand2 add_76_82_g1224 (.a(add_76_82_n_936), .b(add_76_82_n_1097), .y(add_76_82_n_916));
nand2 add_76_82_g1225 (.a(add_76_82_n_938), .b(add_76_82_n_1095), .y(add_76_82_n_918));
nand2 add_76_82_g1226 (.a(add_76_82_n_955), .b(add_76_82_n_1090), .y(add_76_82_n_920));
nor2 add_76_82_g1227 (.a(add_76_82_n_939), .b(n_2577), .y(add_76_82_n_922));
nor2 add_76_82_g1228 (.a(add_76_82_n_937), .b(add_76_82_n_1298), .y(add_76_82_n_923));
nor2 add_76_82_g1231 (.a(add_76_82_n_939), .b(add_76_82_n_1236), .y(add_76_82_n_928));
nand2 add_76_82_g1232 (.a(add_76_82_n_955), .b(add_76_82_n_1058), .y(add_76_82_n_930));
nor2 add_76_82_g1233 (.a(add_76_82_n_956), .b(add_76_82_n_1296), .y(add_76_82_n_931));
nor2 add_76_82_g1235 (.a(add_76_82_n_937), .b(add_76_82_n_1028), .y(add_76_82_n_933));
nand2 add_76_82_g1236 (.a(add_76_82_n_938), .b(add_76_82_n_1057), .y(add_76_82_n_934));
inv add_76_82_g1238 (.a(add_76_82_n_936), .y(add_76_82_n_937));
inv add_76_82_g1239 (.a(add_76_82_n_938), .y(add_76_82_n_939));
nand2 add_76_82_g1240 (.a(add_76_82_n_974), .b(add_76_82_n_1215), .y(add_76_82_n_940));
nand2 add_76_82_g1241 (.a(add_76_82_n_976), .b(add_76_82_n_979), .y(add_76_82_n_941));
nor2 add_76_82_g1242 (.a(add_76_82_n_1010), .b(add_76_82_n_1278), .y(add_76_82_n_944));
nand2 add_76_82_g1243 (.a(add_76_82_n_975), .b(add_76_82_n_1291), .y(add_76_82_n_945));
nor2 add_76_82_g1244 (.a(add_76_82_n_980), .b(add_76_82_n_1299), .y(add_76_82_n_946));
nand2 add_76_82_g1245 (.a(add_76_82_n_1013), .b(add_76_82_n_1228), .y(add_76_82_n_948));
nand2 add_76_82_g1246 (.a(add_76_82_n_979), .b(add_76_82_n_1094), .y(add_76_82_n_949));
nor2 add_76_82_g1247 (.a(add_76_82_n_1007), .b(add_76_82_n_1271), .y(add_76_82_n_951));
nand2 add_76_82_g1249 (.a(add_76_82_n_1009), .b(add_76_82_n_1069), .y(add_76_82_n_954));
nand2 add_76_82_g1250 (.a(add_76_82_n_1012), .b(add_76_82_n_1068), .y(add_76_82_n_936));
nand2 add_76_82_g1251 (.a(add_76_82_n_991), .b(add_76_82_n_1049), .y(add_76_82_n_938));
inv add_76_82_g1252 (.a(add_76_82_n_955), .y(add_76_82_n_956));
nand2 add_76_82_g1254 (.a(add_76_82_n_1000), .b(add_76_82_n_1072), .y(add_76_82_n_959));
nor2 add_76_82_g1255 (.a(add_76_82_n_1015), .b(add_76_82_n_1289), .y(add_76_82_n_960));
nor2 add_76_82_g1256 (.a(add_76_82_n_998), .b(add_76_82_n_1265), .y(add_76_82_n_961));
nor2 add_76_82_g1258 (.a(add_76_82_n_980), .b(add_76_82_n_1030), .y(add_76_82_n_963));
nand2 add_76_82_g1259 (.a(add_76_82_n_1019), .b(add_76_82_n_1073), .y(add_76_82_n_966));
nor2 add_76_82_g1260 (.a(add_76_82_n_980), .b(add_76_82_n_1041), .y(add_76_82_n_967));
nor2 add_76_82_g1261 (.a(add_76_82_n_1004), .b(add_76_82_n_980), .y(add_76_82_n_969));
nor2 add_76_82_g1262 (.a(add_76_82_n_1005), .b(add_76_82_n_980), .y(add_76_82_n_971));
nand2 add_76_82_g1264 (.a(add_76_82_n_1018), .b(add_76_82_n_1048), .y(add_76_82_n_955));
inv add_76_82_g1266 (.a(add_76_82_n_989), .y(add_76_82_n_974));
inv add_76_82_g1267 (.a(add_76_82_n_992), .y(add_76_82_n_975));
inv add_76_82_g1269 (.a(add_76_82_n_979), .y(add_76_82_n_980));
nor2 add_76_82_g1270 (.a(add_76_82_n_1040), .b(add_76_82_n_1298), .y(add_76_82_n_981));
nand2 add_76_82_g1271 (.a(add_76_82_n_1039), .b(add_76_82_n_1097), .y(add_76_82_n_984));
nor2 add_76_82_g1272 (.a(n_2578), .b(add_76_82_n_1236), .y(add_76_82_n_986));
nor2 add_76_82_g1273 (.a(add_76_82_n_1037), .b(add_76_82_n_1300), .y(add_76_82_n_989));
nand2 add_76_82_g1274 (.a(add_76_82_n_1034), .b(add_76_82_n_1084), .y(add_76_82_n_991));
nor2 add_76_82_g1275 (.a(add_76_82_n_1063), .b(add_76_82_n_1233), .y(add_76_82_n_992));
nand2 add_76_82_g1277 (.a(add_76_82_n_1044), .b(add_76_82_n_1095), .y(add_76_82_n_996));
nor2 add_76_82_g1278 (.a(add_76_82_n_1032), .b(add_76_82_n_1203), .y(add_76_82_n_998));
nand2 add_76_82_g1279 (.a(add_76_82_n_1038), .b(add_76_82_n_1082), .y(add_76_82_n_1000));
nor2 add_76_82_g1280 (.a(add_76_82_n_1041), .b(add_76_82_n_1296), .y(add_76_82_n_976));
nor2 add_76_82_g1282 (.a(add_76_82_n_1031), .b(add_76_82_n_1040), .y(add_76_82_n_979));
nor2 add_76_82_g1284 (.a(add_76_82_n_1061), .b(add_76_82_n_1302), .y(add_76_82_n_1007));
nand2 add_76_82_g1285 (.a(add_76_82_n_1060), .b(add_76_82_n_1081), .y(add_76_82_n_1009));
nor2 add_76_82_g1286 (.a(add_76_82_n_1035), .b(add_76_82_n_1230), .y(add_76_82_n_1010));
nand2 add_76_82_g1287 (.a(add_76_82_n_1062), .b(add_76_82_n_1086), .y(add_76_82_n_1012));
nand2 add_76_82_g1288 (.a(add_76_82_n_1034), .b(add_76_82_n_1238), .y(add_76_82_n_1013));
nor2 add_76_82_g1289 (.a(add_76_82_n_1059), .b(add_76_82_n_1231), .y(add_76_82_n_1015));
nand2 add_76_82_g1291 (.a(add_76_82_n_1064), .b(add_76_82_n_1083), .y(add_76_82_n_1018));
nand2 add_76_82_g1292 (.a(add_76_82_n_1036), .b(add_76_82_n_1085), .y(add_76_82_n_1019));
nor2 add_76_82_g1293 (.a(add_76_82_n_1028), .b(add_76_82_n_1040), .y(add_76_82_n_1020));
nand2 add_76_82_g1294 (.a(add_76_82_n_1057), .b(add_76_82_n_1044), .y(add_76_82_n_1022));
nand2 add_76_82_g1295 (.a(add_76_82_n_1058), .b(add_76_82_n_1042), .y(add_76_82_n_1004));
nand2 add_76_82_g1296 (.a(add_76_82_n_1042), .b(add_76_82_n_1090), .y(add_76_82_n_1005));
inv add_76_82_g1298 (.a(add_76_82_n_1035), .y(add_76_82_n_1036));
inv add_76_82_g1299 (.a(add_76_82_n_1037), .y(add_76_82_n_1038));
inv add_76_82_g1300 (.a(add_76_82_n_1040), .y(add_76_82_n_1039));
inv add_76_82_g1301 (.a(add_76_82_n_1041), .y(add_76_82_n_1042));
inv add_76_82_g1302 (.a(n_2578), .y(add_76_82_n_1044));
nor2 add_76_82_g1304 (.a(add_76_82_n_1102), .b(add_76_82_n_1270), .y(add_76_82_n_1048));
nor2 add_76_82_g1305 (.a(add_76_82_n_1104), .b(add_76_82_n_1198), .y(add_76_82_n_1049));
nand2 add_76_82_g1306 (.a(add_76_82_n_1097), .b(add_76_82_n_1301), .y(add_76_82_n_1028));
nand2 add_76_82_g1308 (.a(add_76_82_n_1094), .b(add_76_82_n_1234), .y(add_76_82_n_1030));
nand2 add_76_82_g1309 (.a(add_76_82_n_1082), .b(add_76_82_n_1097), .y(add_76_82_n_1031));
nor2 add_76_82_g1310 (.a(add_76_82_n_1116), .b(add_76_82_n_1258), .y(add_76_82_n_1032));
nand2 add_76_82_g1311 (.a(add_76_82_n_1080), .b(add_76_82_n_1267), .y(add_76_82_n_1034));
nor2 add_76_82_g1312 (.a(add_76_82_n_1122), .b(add_76_82_n_1194), .y(add_76_82_n_1035));
nor2 add_76_82_g1313 (.a(add_76_82_n_1106), .b(add_76_82_n_1261), .y(add_76_82_n_1037));
nand2 add_76_82_g1314 (.a(add_76_82_n_1086), .b(add_76_82_n_1093), .y(add_76_82_n_1040));
nand2 add_76_82_g1315 (.a(add_76_82_n_1083), .b(add_76_82_n_1094), .y(add_76_82_n_1041));
inv add_76_82_g1317 (.a(add_76_82_n_1059), .y(add_76_82_n_1060));
inv add_76_82_g1318 (.a(add_76_82_n_1061), .y(add_76_82_n_1062));
inv add_76_82_g1319 (.a(add_76_82_n_1063), .y(add_76_82_n_1064));
nor2 add_76_82_g1320 (.a(add_76_82_n_1087), .b(add_76_82_n_1231), .y(add_76_82_n_1066));
nor2 add_76_82_g1321 (.a(add_76_82_n_1113), .b(add_76_82_n_1201), .y(add_76_82_n_1068));
nor2 add_76_82_g1322 (.a(add_76_82_n_1111), .b(add_76_82_n_1264), .y(add_76_82_n_1069));
nand2 add_76_82_g1323 (.a(add_76_82_n_1091), .b(add_76_82_n_1238), .y(add_76_82_n_1070));
nor2 add_76_82_g1324 (.a(add_76_82_n_1100), .b(add_76_82_n_1200), .y(add_76_82_n_1072));
nor2 add_76_82_g1325 (.a(add_76_82_n_1112), .b(add_76_82_n_1268), .y(add_76_82_n_1073));
nor2 add_76_82_g1327 (.a(add_76_82_n_1092), .b(add_76_82_n_1302), .y(add_76_82_n_1075));
nor2 add_76_82_g1328 (.a(add_76_82_n_1096), .b(add_76_82_n_1230), .y(add_76_82_n_1057));
nor2 add_76_82_g1329 (.a(add_76_82_n_1089), .b(add_76_82_n_1203), .y(add_76_82_n_1058));
nor2 add_76_82_g1330 (.a(add_76_82_n_1114), .b(add_76_82_n_1257), .y(add_76_82_n_1059));
nor2 add_76_82_g1331 (.a(add_76_82_n_1098), .b(add_76_82_n_1262), .y(add_76_82_n_1061));
nor2 add_76_82_g1332 (.a(add_76_82_n_1117), .b(add_76_82_n_1260), .y(add_76_82_n_1063));
inv add_76_82_g1335 (.a(add_76_82_n_1109), .y(add_76_82_n_1080));
inv add_76_82_g1336 (.a(add_76_82_n_1088), .y(add_76_82_n_1087));
inv add_76_82_g1337 (.a(add_76_82_n_1090), .y(add_76_82_n_1089));
inv add_76_82_g1338 (.a(add_76_82_n_1093), .y(add_76_82_n_1092));
inv add_76_82_g1339 (.a(add_76_82_n_1095), .y(add_76_82_n_1096));
nor2 add_76_82_g1340 (.a(add_76_82_n_1293), .b(add_76_82_n_1275), .y(add_76_82_n_1098));
nor2 add_76_82_g1341 (.a(add_76_82_n_1215), .b(add_76_82_n_1204), .y(add_76_82_n_1100));
nor2 add_76_82_g1342 (.a(add_76_82_n_1291), .b(add_76_82_n_1285), .y(add_76_82_n_1102));
nor2 add_76_82_g1343 (.a(add_76_82_n_1228), .b(add_76_82_n_1295), .y(add_76_82_n_1104));
nor2 add_76_82_g1344 (.a(add_76_82_n_1217), .b(add_76_82_n_1286), .y(add_76_82_n_1106));
nor2 add_76_82_g1346 (.a(add_76_82_n_1276), .b(add_76_82_n_1223), .y(add_76_82_n_1109));
nor2 add_76_82_g1347 (.a(add_76_82_n_1290), .b(add_76_82_n_1224), .y(add_76_82_n_1111));
nor2 add_76_82_g1348 (.a(add_76_82_n_1279), .b(add_76_82_n_1226), .y(add_76_82_n_1112));
nor2 add_76_82_g1349 (.a(add_76_82_n_1272), .b(add_76_82_n_1222), .y(add_76_82_n_1113));
nor2 add_76_82_g1350 (.a(add_76_82_n_1210), .b(add_76_82_n_1273), .y(add_76_82_n_1114));
nor2 add_76_82_g1351 (.a(add_76_82_n_1219), .b(add_76_82_n_1214), .y(add_76_82_n_1116));
nor2 add_76_82_g1352 (.a(add_76_82_n_1212), .b(add_76_82_n_1284), .y(add_76_82_n_1117));
nor2 add_76_82_g1355 (.a(add_76_82_n_1206), .b(add_76_82_n_1277), .y(add_76_82_n_1122));
nor2 add_76_82_g1357 (.a(add_76_82_n_1224), .b(add_76_82_n_1231), .y(add_76_82_n_1081));
nor2 add_76_82_g1358 (.a(add_76_82_n_1204), .b(add_76_82_n_1300), .y(add_76_82_n_1082));
nor2 add_76_82_g1359 (.a(add_76_82_n_1285), .b(add_76_82_n_1233), .y(add_76_82_n_1083));
nor2 add_76_82_g1360 (.a(add_76_82_n_1295), .b(add_76_82_n_1237), .y(add_76_82_n_1084));
nor2 add_76_82_g1361 (.a(add_76_82_n_1226), .b(add_76_82_n_1230), .y(add_76_82_n_1085));
nor2 add_76_82_g1362 (.a(add_76_82_n_1222), .b(add_76_82_n_1302), .y(add_76_82_n_1086));
nor2 add_76_82_g1363 (.a(add_76_82_n_1273), .b(n_1843), .y(add_76_82_n_1088));
nor2 add_76_82_g1364 (.a(add_76_82_n_1214), .b(add_76_82_n_1296), .y(add_76_82_n_1090));
nor2 add_76_82_g1365 (.a(add_76_82_n_1223), .b(add_76_82_n_1208), .y(add_76_82_n_1091));
nor2 add_76_82_g1366 (.a(add_76_82_n_1275), .b(add_76_82_n_1232), .y(add_76_82_n_1093));
nor2 add_76_82_g1367 (.a(add_76_82_n_1284), .b(add_76_82_n_1299), .y(add_76_82_n_1094));
nor2 add_76_82_g1368 (.a(add_76_82_n_1277), .b(add_76_82_n_1236), .y(add_76_82_n_1095));
nor2 add_76_82_g1369 (.a(add_76_82_n_1286), .b(add_76_82_n_1298), .y(add_76_82_n_1097));
xor2 add_76_82_g1370 (.a(n_688), .b(sum_0_), .y(n_849));
nor2 add_76_82_g1372 (.a(add_76_82_n_1209), .b(n_1843), .y(add_76_82_n_1144));
nand2 add_76_82_g1374 (.a(add_76_82_n_1276), .b(add_76_82_n_1207), .y(add_76_82_n_1148));
nor2 add_76_82_g1377 (.a(add_76_82_n_1265), .b(add_76_82_n_1203), .y(add_76_82_n_1153));
nor2 add_76_82_g1385 (.a(add_76_82_n_1292), .b(add_76_82_n_1232), .y(add_76_82_n_1168));
xor2 add_76_82_g1399 (.a(n_719), .b(sum_31_), .y(add_76_82_n_1191));
inv add_76_82_g1401 (.a(add_76_82_n_1239), .y(add_76_82_n_1194));
inv add_76_82_g1402 (.a(n_1866), .y(add_76_82_n_1196));
inv add_76_82_g1403 (.a(add_76_82_n_1199), .y(add_76_82_n_1198));
inv add_76_82_g1404 (.a(add_76_82_n_1242), .y(add_76_82_n_1200));
inv add_76_82_g1405 (.a(add_76_82_n_1243), .y(add_76_82_n_1201));
inv add_76_82_g1407 (.a(add_76_82_n_1206), .y(add_76_82_n_1205));
inv add_76_82_g1408 (.a(add_76_82_n_1208), .y(add_76_82_n_1207));
inv add_76_82_g1409 (.a(add_76_82_n_1210), .y(add_76_82_n_1209));
inv add_76_82_g1410 (.a(add_76_82_n_1212), .y(add_76_82_n_1211));
inv add_76_82_g1411 (.a(add_76_82_n_1214), .y(add_76_82_n_1213));
inv add_76_82_g1412 (.a(add_76_82_n_1217), .y(add_76_82_n_1216));
inv add_76_82_g1413 (.a(add_76_82_n_1219), .y(add_76_82_n_1218));
inv add_76_82_g1414 (.a(add_76_82_n_1226), .y(add_76_82_n_1225));
inv add_76_82_g1415 (.a(add_76_82_n_1228), .y(add_76_82_n_1227));
inv add_76_82_g1416 (.a(add_76_82_n_1230), .y(add_76_82_n_1229));
inv add_76_82_g1417 (.a(add_76_82_n_1233), .y(add_76_82_n_1234));
inv add_76_82_g1418 (.a(add_76_82_n_1236), .y(add_76_82_n_1235));
inv add_76_82_g1419 (.a(add_76_82_n_1237), .y(add_76_82_n_1238));
nand2 add_76_82_g1420 (.a(n_701), .b(sum_13_), .y(add_76_82_n_1239));
nand2 add_76_82_g1423 (.a(n_699), .b(sum_11_), .y(add_76_82_n_1199));
nand2 add_76_82_g1424 (.a(n_711), .b(sum_23_), .y(add_76_82_n_1242));
nand2 add_76_82_g1425 (.a(n_707), .b(sum_19_), .y(add_76_82_n_1243));
nor2 add_76_82_g1427 (.a(n_718), .b(sum_30_), .y(add_76_82_n_1203));
nor2 add_76_82_g1428 (.a(n_711), .b(sum_23_), .y(add_76_82_n_1204));
nand2 add_76_82_g1429 (.a(n_700), .b(sum_12_), .y(add_76_82_n_1206));
nor2 add_76_82_g1430 (.a(n_696), .b(sum_8_), .y(add_76_82_n_1208));
nand2 add_76_82_g1431 (.a(n_1842), .b(sum_4_), .y(add_76_82_n_1210));
nand2 add_76_82_g1432 (.a(n_712), .b(sum_24_), .y(add_76_82_n_1212));
nor2 add_76_82_g1433 (.a(n_717), .b(sum_29_), .y(add_76_82_n_1214));
nand2 add_76_82_g1434 (.a(n_710), .b(sum_22_), .y(add_76_82_n_1215));
nand2 add_76_82_g1435 (.a(n_708), .b(sum_20_), .y(add_76_82_n_1217));
nand2 add_76_82_g1436 (.a(n_716), .b(sum_28_), .y(add_76_82_n_1219));
nor2 add_76_82_g1439 (.a(n_707), .b(sum_19_), .y(add_76_82_n_1222));
nor2 add_76_82_g1440 (.a(n_697), .b(sum_9_), .y(add_76_82_n_1223));
nor2 add_76_82_g1441 (.a(n_695), .b(sum_7_), .y(add_76_82_n_1224));
nor2 add_76_82_g1442 (.a(n_703), .b(sum_15_), .y(add_76_82_n_1226));
nand2 add_76_82_g1443 (.a(n_698), .b(sum_10_), .y(add_76_82_n_1228));
nor2 add_76_82_g1444 (.a(n_702), .b(sum_14_), .y(add_76_82_n_1230));
nor2 add_76_82_g1445 (.a(n_694), .b(sum_6_), .y(add_76_82_n_1231));
nor2 add_76_82_g1446 (.a(n_704), .b(sum_16_), .y(add_76_82_n_1232));
nor2 add_76_82_g1447 (.a(n_714), .b(sum_26_), .y(add_76_82_n_1233));
nor2 add_76_82_g1448 (.a(n_700), .b(sum_12_), .y(add_76_82_n_1236));
nor2 add_76_82_g1449 (.a(n_698), .b(sum_10_), .y(add_76_82_n_1237));
inv add_76_82_g1450 (.a(add_76_82_n_1303), .y(add_76_82_n_1257));
inv add_76_82_g1451 (.a(add_76_82_n_1259), .y(add_76_82_n_1258));
inv add_76_82_g1452 (.a(add_76_82_n_1306), .y(add_76_82_n_1260));
inv add_76_82_g1453 (.a(add_76_82_n_1307), .y(add_76_82_n_1261));
inv add_76_82_g1454 (.a(add_76_82_n_1263), .y(add_76_82_n_1262));
inv add_76_82_g1455 (.a(add_76_82_n_1308), .y(add_76_82_n_1264));
inv add_76_82_g1456 (.a(add_76_82_n_1311), .y(add_76_82_n_1265));
inv add_76_82_g1457 (.a(add_76_82_n_1267), .y(add_76_82_n_1266));
inv add_76_82_g1458 (.a(add_76_82_n_1269), .y(add_76_82_n_1268));
inv add_76_82_g1459 (.a(add_76_82_n_1318), .y(add_76_82_n_1270));
inv add_76_82_g1460 (.a(add_76_82_n_1272), .y(add_76_82_n_1271));
inv add_76_82_g1461 (.a(add_76_82_n_1275), .y(add_76_82_n_1274));
inv add_76_82_g1462 (.a(add_76_82_n_1279), .y(add_76_82_n_1278));
inv add_76_82_g1465 (.a(n_2901), .y(add_76_82_n_1287));
inv add_76_82_g1466 (.a(add_76_82_n_1290), .y(add_76_82_n_1289));
inv add_76_82_g1467 (.a(add_76_82_n_1293), .y(add_76_82_n_1292));
inv add_76_82_g1468 (.a(add_76_82_n_1295), .y(add_76_82_n_1294));
inv add_76_82_g1469 (.a(add_76_82_n_1298), .y(add_76_82_n_1297));
inv add_76_82_g1470 (.a(add_76_82_n_1300), .y(add_76_82_n_1301));
nand2 add_76_82_g1471 (.a(n_693), .b(sum_5_), .y(add_76_82_n_1303));
nand2 add_76_82_g1472 (.a(n_717), .b(sum_29_), .y(add_76_82_n_1259));
nand2 add_76_82_g1473 (.a(n_713), .b(sum_25_), .y(add_76_82_n_1306));
nand2 add_76_82_g1474 (.a(n_709), .b(sum_21_), .y(add_76_82_n_1307));
nand2 add_76_82_g1475 (.a(n_705), .b(sum_17_), .y(add_76_82_n_1263));
nand2 add_76_82_g1476 (.a(n_695), .b(sum_7_), .y(add_76_82_n_1308));
nand2 add_76_82_g1477 (.a(n_718), .b(sum_30_), .y(add_76_82_n_1311));
nand2 add_76_82_g1478 (.a(n_697), .b(sum_9_), .y(add_76_82_n_1267));
nand2 add_76_82_g1479 (.a(n_703), .b(sum_15_), .y(add_76_82_n_1269));
nand2 add_76_82_g1480 (.a(n_715), .b(sum_27_), .y(add_76_82_n_1318));
nand2 add_76_82_g1481 (.a(n_706), .b(sum_18_), .y(add_76_82_n_1272));
nor2 add_76_82_g1482 (.a(n_693), .b(sum_5_), .y(add_76_82_n_1273));
nor2 add_76_82_g1483 (.a(n_705), .b(sum_17_), .y(add_76_82_n_1275));
nand2 add_76_82_g1484 (.a(n_696), .b(sum_8_), .y(add_76_82_n_1276));
nor2 add_76_82_g1485 (.a(n_701), .b(sum_13_), .y(add_76_82_n_1277));
nand2 add_76_82_g1486 (.a(n_702), .b(sum_14_), .y(add_76_82_n_1279));
nor2 add_76_82_g1489 (.a(n_713), .b(sum_25_), .y(add_76_82_n_1284));
nor2 add_76_82_g1490 (.a(n_715), .b(sum_27_), .y(add_76_82_n_1285));
nor2 add_76_82_g1491 (.a(n_709), .b(sum_21_), .y(add_76_82_n_1286));
nand2 add_76_82_g1493 (.a(n_694), .b(sum_6_), .y(add_76_82_n_1290));
nand2 add_76_82_g1494 (.a(n_714), .b(sum_26_), .y(add_76_82_n_1291));
nand2 add_76_82_g1495 (.a(n_704), .b(sum_16_), .y(add_76_82_n_1293));
nor2 add_76_82_g1496 (.a(n_699), .b(sum_11_), .y(add_76_82_n_1295));
nor2 add_76_82_g1497 (.a(n_716), .b(sum_28_), .y(add_76_82_n_1296));
nor2 add_76_82_g1498 (.a(n_708), .b(sum_20_), .y(add_76_82_n_1298));
nor2 add_76_82_g1499 (.a(n_712), .b(sum_24_), .y(add_76_82_n_1299));
nor2 add_76_82_g1500 (.a(n_710), .b(sum_22_), .y(add_76_82_n_1300));
nor2 add_76_82_g1501 (.a(n_706), .b(sum_18_), .y(add_76_82_n_1302));
xor2 add_76_69_g942 (.a(add_76_69_n_625), .b(add_76_69_n_981), .y(n_940));
xor2 add_76_69_g950 (.a(add_76_69_n_631), .b(add_76_69_n_994), .y(n_943));
nand2 add_76_69_g953 (.a(add_76_69_n_668), .b(add_76_69_n_660), .y(add_76_69_n_625));
nand2 add_76_69_g959 (.a(add_76_69_n_666), .b(add_76_69_n_653), .y(add_76_69_n_631));
nor2 add_76_69_g978 (.a(add_76_69_n_664), .b(add_76_69_n_750), .y(add_76_69_n_651));
nand2 add_76_69_g979 (.a(n_3843), .b(add_76_69_n_772), .y(add_76_69_n_653));
nand2 add_76_69_g980 (.a(n_3843), .b(add_76_69_n_788), .y(add_76_69_n_654));
nand2 add_76_69_g981 (.a(n_3843), .b(add_76_69_n_768), .y(add_76_69_n_655));
nand2 add_76_69_g982 (.a(n_3843), .b(add_76_69_n_781), .y(add_76_69_n_656));
nor2 add_76_69_g984 (.a(add_76_69_n_664), .b(add_76_69_n_842), .y(add_76_69_n_658));
nand2 add_76_69_g985 (.a(n_3843), .b(add_76_69_n_823), .y(add_76_69_n_659));
nand2 add_76_69_g986 (.a(n_3843), .b(add_76_69_n_774), .y(add_76_69_n_660));
nand2 add_76_69_g987 (.a(n_3843), .b(add_76_69_n_776), .y(add_76_69_n_661));
inv add_76_69_g989 (.a(n_3843), .y(add_76_69_n_664));
nand2 add_76_69_g990 (.a(add_76_69_n_684), .b(add_76_69_n_716), .y(add_76_69_n_665));
nor2 add_76_69_g991 (.a(add_76_69_n_700), .b(add_76_69_n_709), .y(add_76_69_n_666));
nor2 add_76_69_g993 (.a(add_76_69_n_699), .b(add_76_69_n_715), .y(add_76_69_n_668));
nor2 add_76_69_g994 (.a(add_76_69_n_696), .b(add_76_69_n_761), .y(add_76_69_n_669));
nor2 add_76_69_g1000 (.a(add_76_69_n_701), .b(add_76_69_n_763), .y(add_76_69_n_674));
xor2 add_76_69_g1001 (.a(add_76_69_n_705), .b(add_76_69_n_988), .y(n_874));
inv add_76_69_g1009 (.a(add_76_69_n_685), .y(add_76_69_n_683));
nand2 add_76_69_g1010 (.a(n_2321), .b(add_76_69_n_780), .y(add_76_69_n_684));
nor2 add_76_69_g1011 (.a(add_76_69_n_705), .b(add_76_69_n_1034), .y(add_76_69_n_685));
nand2 add_76_69_g1014 (.a(add_76_69_n_706), .b(add_76_69_n_783), .y(add_76_69_n_690));
nand2 add_76_69_g1015 (.a(add_76_69_n_706), .b(add_76_69_n_897), .y(add_76_69_n_692));
nor2 add_76_69_g1018 (.a(n_2320), .b(add_76_69_n_843), .y(add_76_69_n_696));
nor2 add_76_69_g1019 (.a(add_76_69_n_705), .b(add_76_69_n_795), .y(add_76_69_n_697));
nor2 add_76_69_g1020 (.a(add_76_69_n_705), .b(add_76_69_n_845), .y(add_76_69_n_698));
nor2 add_76_69_g1021 (.a(n_2320), .b(add_76_69_n_807), .y(add_76_69_n_699));
nor2 add_76_69_g1022 (.a(n_2320), .b(add_76_69_n_806), .y(add_76_69_n_700));
nor2 add_76_69_g1023 (.a(n_2320), .b(add_76_69_n_861), .y(add_76_69_n_701));
inv add_76_69_g1026 (.a(add_76_69_n_705), .y(add_76_69_n_706));
nand2 add_76_69_g1027 (.a(add_76_69_n_732), .b(add_76_69_n_863), .y(add_76_69_n_707));
nand2 add_76_69_g1029 (.a(add_76_69_n_736), .b(add_76_69_n_765), .y(add_76_69_n_709));
nand2 add_76_69_g1030 (.a(add_76_69_n_723), .b(add_76_69_n_867), .y(add_76_69_n_710));
nor2 add_76_69_g1031 (.a(add_76_69_n_722), .b(add_76_69_n_1092), .y(add_76_69_n_711));
nor2 add_76_69_g1034 (.a(add_76_69_n_760), .b(add_76_69_n_735), .y(add_76_69_n_705));
nor2 add_76_69_g1036 (.a(add_76_69_n_738), .b(add_76_69_n_1016), .y(add_76_69_n_714));
nand2 add_76_69_g1037 (.a(add_76_69_n_727), .b(add_76_69_n_832), .y(add_76_69_n_715));
nor2 add_76_69_g1038 (.a(add_76_69_n_737), .b(add_76_69_n_1099), .y(add_76_69_n_716));
nor2 add_76_69_g1039 (.a(add_76_69_n_740), .b(add_76_69_n_756), .y(add_76_69_n_717));
nor2 add_76_69_g1044 (.a(add_76_69_n_744), .b(add_76_69_n_1042), .y(add_76_69_n_722));
nand2 add_76_69_g1045 (.a(add_76_69_n_745), .b(add_76_69_n_898), .y(add_76_69_n_723));
nand2 add_76_69_g1047 (.a(add_76_69_n_761), .b(add_76_69_n_894), .y(add_76_69_n_727));
nor2 add_76_69_g1048 (.a(add_76_69_n_746), .b(add_76_69_n_831), .y(add_76_69_n_729));
nand2 add_76_69_g1050 (.a(add_76_69_n_743), .b(add_76_69_n_900), .y(add_76_69_n_732));
nand2 add_76_69_g1051 (.a(n_2927), .b(add_76_69_n_1022), .y(add_76_69_n_734));
nor2 add_76_69_g1052 (.a(add_76_69_n_748), .b(n_2944), .y(add_76_69_n_735));
nand2 add_76_69_g1053 (.a(add_76_69_n_761), .b(add_76_69_n_862), .y(add_76_69_n_736));
nor2 add_76_69_g1054 (.a(add_76_69_n_762), .b(add_76_69_n_1105), .y(add_76_69_n_737));
nor2 add_76_69_g1055 (.a(add_76_69_n_746), .b(add_76_69_n_1107), .y(add_76_69_n_738));
nor2 add_76_69_g1056 (.a(add_76_69_n_744), .b(add_76_69_n_834), .y(add_76_69_n_740));
nand2 add_76_69_g1057 (.a(add_76_69_n_745), .b(add_76_69_n_860), .y(add_76_69_n_741));
nand2 add_76_69_g1058 (.a(n_2927), .b(add_76_69_n_870), .y(add_76_69_n_742));
inv add_76_69_g1059 (.a(add_76_69_n_743), .y(add_76_69_n_744));
inv add_76_69_g1060 (.a(add_76_69_n_745), .y(add_76_69_n_746));
inv add_76_69_g1061 (.a(n_2927), .y(add_76_69_n_748));
nor2 add_76_69_g1062 (.a(add_76_69_n_791), .b(add_76_69_n_1024), .y(add_76_69_n_749));
nand2 add_76_69_g1063 (.a(add_76_69_n_780), .b(add_76_69_n_781), .y(add_76_69_n_750));
nor2 add_76_69_g1064 (.a(add_76_69_n_782), .b(add_76_69_n_1043), .y(add_76_69_n_753));
nand2 add_76_69_g1065 (.a(add_76_69_n_813), .b(add_76_69_n_1095), .y(add_76_69_n_755));
nand2 add_76_69_g1066 (.a(add_76_69_n_779), .b(add_76_69_n_1018), .y(add_76_69_n_756));
nand2 add_76_69_g1067 (.a(add_76_69_n_781), .b(add_76_69_n_901), .y(add_76_69_n_757));
nor2 add_76_69_g1068 (.a(add_76_69_n_810), .b(add_76_69_n_1097), .y(add_76_69_n_759));
nand2 add_76_69_g1069 (.a(add_76_69_n_809), .b(add_76_69_n_877), .y(add_76_69_n_760));
nand2 add_76_69_g1070 (.a(add_76_69_n_812), .b(add_76_69_n_851), .y(add_76_69_n_743));
nand2 add_76_69_g1071 (.a(add_76_69_n_799), .b(add_76_69_n_852), .y(add_76_69_n_745));
inv add_76_69_g1073 (.a(add_76_69_n_761), .y(add_76_69_n_762));
nand2 add_76_69_g1074 (.a(add_76_69_n_821), .b(add_76_69_n_1085), .y(add_76_69_n_763));
nor2 add_76_69_g1076 (.a(add_76_69_n_802), .b(add_76_69_n_1071), .y(add_76_69_n_765));
nand2 add_76_69_g1077 (.a(add_76_69_n_820), .b(add_76_69_n_879), .y(add_76_69_n_766));
nand2 add_76_69_g1078 (.a(add_76_69_n_794), .b(add_76_69_n_878), .y(add_76_69_n_767));
nor2 add_76_69_g1079 (.a(add_76_69_n_782), .b(add_76_69_n_861), .y(add_76_69_n_768));
nor2 add_76_69_g1080 (.a(n_2943), .b(add_76_69_n_1080), .y(add_76_69_n_771));
nor2 add_76_69_g1081 (.a(add_76_69_n_806), .b(add_76_69_n_782), .y(add_76_69_n_772));
nor2 add_76_69_g1082 (.a(add_76_69_n_807), .b(add_76_69_n_782), .y(add_76_69_n_774));
nor2 add_76_69_g1083 (.a(add_76_69_n_782), .b(add_76_69_n_843), .y(add_76_69_n_776));
nand2 add_76_69_g1084 (.a(add_76_69_n_819), .b(add_76_69_n_1032), .y(add_76_69_n_778));
nand2 add_76_69_g1085 (.a(add_76_69_n_793), .b(add_76_69_n_847), .y(add_76_69_n_761));
inv add_76_69_g1086 (.a(add_76_69_n_797), .y(add_76_69_n_779));
inv add_76_69_g1087 (.a(add_76_69_n_781), .y(add_76_69_n_782));
nor2 add_76_69_g1088 (.a(add_76_69_n_845), .b(add_76_69_n_1107), .y(add_76_69_n_783));
nor2 add_76_69_g1089 (.a(add_76_69_n_831), .b(add_76_69_n_845), .y(add_76_69_n_786));
nor2 add_76_69_g1090 (.a(add_76_69_n_842), .b(add_76_69_n_1042), .y(add_76_69_n_788));
nor2 add_76_69_g1091 (.a(add_76_69_n_835), .b(add_76_69_n_1104), .y(add_76_69_n_791));
nand2 add_76_69_g1092 (.a(add_76_69_n_838), .b(add_76_69_n_887), .y(add_76_69_n_793));
nand2 add_76_69_g1093 (.a(add_76_69_n_864), .b(add_76_69_n_886), .y(add_76_69_n_794));
nand2 add_76_69_g1094 (.a(add_76_69_n_846), .b(add_76_69_n_898), .y(add_76_69_n_795));
nor2 add_76_69_g1095 (.a(add_76_69_n_863), .b(add_76_69_n_1108), .y(add_76_69_n_797));
nand2 add_76_69_g1096 (.a(add_76_69_n_840), .b(add_76_69_n_888), .y(add_76_69_n_799));
nand2 add_76_69_g1097 (.a(add_76_69_n_841), .b(add_76_69_n_900), .y(add_76_69_n_800));
nor2 add_76_69_g1098 (.a(add_76_69_n_832), .b(add_76_69_n_1084), .y(add_76_69_n_802));
nor2 add_76_69_g1099 (.a(add_76_69_n_843), .b(add_76_69_n_1105), .y(add_76_69_n_780));
nor2 add_76_69_g1100 (.a(add_76_69_n_833), .b(add_76_69_n_842), .y(add_76_69_n_781));
nand2 add_76_69_g1102 (.a(n_2942), .b(add_76_69_n_890), .y(add_76_69_n_809));
nor2 add_76_69_g1103 (.a(add_76_69_n_867), .b(add_76_69_n_1103), .y(add_76_69_n_810));
nand2 add_76_69_g1104 (.a(add_76_69_n_836), .b(add_76_69_n_885), .y(add_76_69_n_812));
nand2 add_76_69_g1105 (.a(add_76_69_n_840), .b(add_76_69_n_1040), .y(add_76_69_n_813));
nand2 add_76_69_g1106 (.a(add_76_69_n_869), .b(add_76_69_n_908), .y(add_76_69_n_815));
nand2 add_76_69_g1108 (.a(add_76_69_n_869), .b(add_76_69_n_1014), .y(add_76_69_n_819));
nand2 add_76_69_g1109 (.a(add_76_69_n_868), .b(add_76_69_n_889), .y(add_76_69_n_820));
nand2 add_76_69_g1110 (.a(add_76_69_n_838), .b(add_76_69_n_1037), .y(add_76_69_n_821));
nor2 add_76_69_g1111 (.a(add_76_69_n_834), .b(add_76_69_n_842), .y(add_76_69_n_823));
nand2 add_76_69_g1112 (.a(add_76_69_n_860), .b(add_76_69_n_846), .y(add_76_69_n_825));
nand2 add_76_69_g1113 (.a(add_76_69_n_844), .b(add_76_69_n_862), .y(add_76_69_n_806));
nand2 add_76_69_g1114 (.a(add_76_69_n_844), .b(add_76_69_n_894), .y(add_76_69_n_807));
inv add_76_69_g1116 (.a(add_76_69_n_838), .y(add_76_69_n_837));
inv add_76_69_g1117 (.a(add_76_69_n_840), .y(add_76_69_n_839));
inv add_76_69_g1118 (.a(add_76_69_n_842), .y(add_76_69_n_841));
inv add_76_69_g1119 (.a(add_76_69_n_843), .y(add_76_69_n_844));
inv add_76_69_g1120 (.a(add_76_69_n_845), .y(add_76_69_n_846));
nor2 add_76_69_g1121 (.a(add_76_69_n_903), .b(add_76_69_n_1004), .y(add_76_69_n_847));
nor2 add_76_69_g1123 (.a(add_76_69_n_918), .b(add_76_69_n_998), .y(add_76_69_n_851));
nor2 add_76_69_g1124 (.a(add_76_69_n_905), .b(add_76_69_n_1002), .y(add_76_69_n_852));
nand2 add_76_69_g1125 (.a(add_76_69_n_889), .b(add_76_69_n_898), .y(add_76_69_n_831));
nor2 add_76_69_g1126 (.a(add_76_69_n_912), .b(add_76_69_n_1011), .y(add_76_69_n_832));
nand2 add_76_69_g1127 (.a(add_76_69_n_886), .b(add_76_69_n_900), .y(add_76_69_n_833));
nand2 add_76_69_g1128 (.a(add_76_69_n_900), .b(add_76_69_n_1109), .y(add_76_69_n_834));
nor2 add_76_69_g1129 (.a(add_76_69_n_921), .b(add_76_69_n_1066), .y(add_76_69_n_835));
nand2 add_76_69_g1130 (.a(add_76_69_n_909), .b(add_76_69_n_1009), .y(add_76_69_n_838));
nand2 add_76_69_g1131 (.a(add_76_69_n_883), .b(add_76_69_n_1007), .y(add_76_69_n_840));
nand2 add_76_69_g1132 (.a(add_76_69_n_885), .b(add_76_69_n_896), .y(add_76_69_n_842));
nand2 add_76_69_g1133 (.a(add_76_69_n_901), .b(add_76_69_n_887), .y(add_76_69_n_843));
nand2 add_76_69_g1134 (.a(add_76_69_n_888), .b(add_76_69_n_897), .y(add_76_69_n_845));
inv add_76_69_g1135 (.a(add_76_69_n_863), .y(add_76_69_n_864));
inv add_76_69_g1137 (.a(add_76_69_n_867), .y(add_76_69_n_868));
nor2 add_76_69_g1138 (.a(n_2945), .b(add_76_69_n_1101), .y(add_76_69_n_870));
nand2 add_76_69_g1139 (.a(add_76_69_n_897), .b(add_76_69_n_1040), .y(add_76_69_n_872));
nor2 add_76_69_g1140 (.a(add_76_69_n_915), .b(add_76_69_n_1005), .y(add_76_69_n_874));
nor2 add_76_69_g1141 (.a(add_76_69_n_895), .b(add_76_69_n_1104), .y(add_76_69_n_875));
nor2 add_76_69_g1142 (.a(add_76_69_n_911), .b(add_76_69_n_1068), .y(add_76_69_n_877));
nor2 add_76_69_g1143 (.a(add_76_69_n_925), .b(add_76_69_n_999), .y(add_76_69_n_878));
nor2 add_76_69_g1144 (.a(add_76_69_n_902), .b(add_76_69_n_1069), .y(add_76_69_n_879));
nor2 add_76_69_g1145 (.a(add_76_69_n_899), .b(add_76_69_n_1103), .y(add_76_69_n_860));
nand2 add_76_69_g1146 (.a(add_76_69_n_901), .b(add_76_69_n_1037), .y(add_76_69_n_861));
nor2 add_76_69_g1147 (.a(add_76_69_n_893), .b(add_76_69_n_1084), .y(add_76_69_n_862));
nor2 add_76_69_g1148 (.a(add_76_69_n_907), .b(add_76_69_n_1072), .y(add_76_69_n_863));
nor2 add_76_69_g1150 (.a(add_76_69_n_927), .b(add_76_69_n_1067), .y(add_76_69_n_867));
nand2 add_76_69_g1151 (.a(add_76_69_n_884), .b(add_76_69_n_1010), .y(add_76_69_n_869));
inv add_76_69_g1152 (.a(add_76_69_n_919), .y(add_76_69_n_883));
inv add_76_69_g1153 (.a(add_76_69_n_923), .y(add_76_69_n_884));
inv add_76_69_g1155 (.a(add_76_69_n_894), .y(add_76_69_n_893));
inv add_76_69_g1156 (.a(add_76_69_n_896), .y(add_76_69_n_895));
inv add_76_69_g1157 (.a(add_76_69_n_898), .y(add_76_69_n_899));
nor2 add_76_69_g1158 (.a(add_76_69_n_1098), .b(add_76_69_n_1030), .y(add_76_69_n_902));
nor2 add_76_69_g1159 (.a(add_76_69_n_1085), .b(add_76_69_n_1096), .y(add_76_69_n_903));
nor2 add_76_69_g1160 (.a(add_76_69_n_1095), .b(add_76_69_n_1087), .y(add_76_69_n_905));
nor2 add_76_69_g1161 (.a(add_76_69_n_1093), .b(add_76_69_n_1019), .y(add_76_69_n_907));
nor2 add_76_69_g1162 (.a(add_76_69_n_1074), .b(add_76_69_n_1015), .y(add_76_69_n_908));
nand2 add_76_69_g1163 (.a(add_76_69_n_1027), .b(add_76_69_n_1076), .y(add_76_69_n_909));
nor2 add_76_69_g1164 (.a(add_76_69_n_1081), .b(add_76_69_n_1091), .y(add_76_69_n_911));
nor2 add_76_69_g1165 (.a(add_76_69_n_1100), .b(add_76_69_n_1083), .y(add_76_69_n_912));
nor2 add_76_69_g1166 (.a(add_76_69_n_1021), .b(add_76_69_n_1078), .y(add_76_69_n_913));
nor2 add_76_69_g1167 (.a(add_76_69_n_1032), .b(add_76_69_n_1074), .y(add_76_69_n_915));
nor2 add_76_69_g1168 (.a(add_76_69_n_1025), .b(add_76_69_n_1026), .y(add_76_69_n_918));
nor2 add_76_69_g1169 (.a(add_76_69_n_1088), .b(add_76_69_n_1079), .y(add_76_69_n_919));
nor2 add_76_69_g1170 (.a(add_76_69_n_1036), .b(add_76_69_n_1077), .y(add_76_69_n_921));
nor2 add_76_69_g1171 (.a(add_76_69_n_1013), .b(add_76_69_n_1001), .y(add_76_69_n_923));
nor2 add_76_69_g1172 (.a(add_76_69_n_1018), .b(add_76_69_n_1073), .y(add_76_69_n_925));
nor2 add_76_69_g1173 (.a(add_76_69_n_1017), .b(add_76_69_n_1028), .y(add_76_69_n_927));
nor2 add_76_69_g1174 (.a(add_76_69_n_1026), .b(add_76_69_n_1104), .y(add_76_69_n_885));
nor2 add_76_69_g1175 (.a(add_76_69_n_1073), .b(add_76_69_n_1108), .y(add_76_69_n_886));
nor2 add_76_69_g1176 (.a(add_76_69_n_1038), .b(add_76_69_n_1096), .y(add_76_69_n_887));
nor2 add_76_69_g1177 (.a(add_76_69_n_1087), .b(add_76_69_n_1039), .y(add_76_69_n_888));
nor2 add_76_69_g1178 (.a(add_76_69_n_1030), .b(add_76_69_n_1103), .y(add_76_69_n_889));
nor2 add_76_69_g1179 (.a(add_76_69_n_1091), .b(add_76_69_n_1101), .y(add_76_69_n_890));
nand2 add_76_69_g1180 (.a(add_76_69_n_1085), .b(add_76_69_n_1037), .y(add_76_69_n_935));
nor2 add_76_69_g1182 (.a(add_76_69_n_1083), .b(add_76_69_n_1105), .y(add_76_69_n_894));
nor2 add_76_69_g1183 (.a(add_76_69_n_1077), .b(add_76_69_n_1090), .y(add_76_69_n_896));
nor2 add_76_69_g1184 (.a(add_76_69_n_1079), .b(add_76_69_n_1034), .y(add_76_69_n_897));
nor2 add_76_69_g1185 (.a(add_76_69_n_1028), .b(add_76_69_n_1107), .y(add_76_69_n_898));
nor2 add_76_69_g1186 (.a(add_76_69_n_1019), .b(add_76_69_n_1042), .y(add_76_69_n_900));
nor2 add_76_69_g1187 (.a(add_76_69_n_1075), .b(add_76_69_n_1043), .y(add_76_69_n_901));
xor2 add_76_69_g1188 (.a(v1_5_), .b(v1_0_), .y(n_850));
nand2 add_76_69_g1191 (.a(add_76_69_n_1018), .b(add_76_69_n_1109), .y(add_76_69_n_948));
nor2 add_76_69_g1193 (.a(add_76_69_n_1031), .b(add_76_69_n_1015), .y(add_76_69_n_952));
nor2 add_76_69_g1194 (.a(add_76_69_n_1005), .b(add_76_69_n_1074), .y(add_76_69_n_954));
nor2 add_76_69_g1199 (.a(add_76_69_n_1035), .b(add_76_69_n_1090), .y(add_76_69_n_964));
nor2 add_76_69_g1207 (.a(add_76_69_n_1080), .b(add_76_69_n_1101), .y(add_76_69_n_977));
nor2 add_76_69_g1209 (.a(add_76_69_n_1071), .b(add_76_69_n_1084), .y(add_76_69_n_981));
nand2 add_76_69_g1210 (.a(add_76_69_n_1010), .b(add_76_69_n_1000), .y(add_76_69_n_983));
nand2 add_76_69_g1213 (.a(add_76_69_n_1088), .b(add_76_69_n_1033), .y(add_76_69_n_988));
xor2 add_76_69_g1217 (.a(v1_31_), .b(v1_27_), .y(add_76_69_n_994));
nor2 add_76_69_g1218 (.a(add_76_69_n_1020), .b(add_76_69_n_1023), .y(add_76_69_n_995));
inv add_76_69_g1219 (.a(add_76_69_n_1044), .y(add_76_69_n_997));
inv add_76_69_g1220 (.a(add_76_69_n_1046), .y(add_76_69_n_998));
inv add_76_69_g1221 (.a(add_76_69_n_1047), .y(add_76_69_n_999));
inv add_76_69_g1222 (.a(add_76_69_n_1001), .y(add_76_69_n_1000));
inv add_76_69_g1223 (.a(add_76_69_n_1003), .y(add_76_69_n_1002));
inv add_76_69_g1224 (.a(add_76_69_n_1048), .y(add_76_69_n_1004));
inv add_76_69_g1225 (.a(add_76_69_n_1051), .y(add_76_69_n_1005));
inv add_76_69_g1226 (.a(add_76_69_n_1007), .y(add_76_69_n_1006));
inv add_76_69_g1227 (.a(add_76_69_n_1009), .y(add_76_69_n_1008));
inv add_76_69_g1228 (.a(add_76_69_n_1012), .y(add_76_69_n_1011));
inv add_76_69_g1229 (.a(add_76_69_n_1015), .y(add_76_69_n_1014));
inv add_76_69_g1230 (.a(add_76_69_n_1017), .y(add_76_69_n_1016));
inv add_76_69_g1231 (.a(add_76_69_n_1021), .y(add_76_69_n_1020));
inv add_76_69_g1232 (.a(add_76_69_n_1023), .y(add_76_69_n_1022));
inv add_76_69_g1233 (.a(add_76_69_n_1025), .y(add_76_69_n_1024));
inv add_76_69_g1234 (.a(add_76_69_n_1060), .y(add_76_69_n_1027));
inv add_76_69_g1235 (.a(add_76_69_n_1030), .y(add_76_69_n_1029));
inv add_76_69_g1236 (.a(add_76_69_n_1032), .y(add_76_69_n_1031));
inv add_76_69_g1237 (.a(add_76_69_n_1034), .y(add_76_69_n_1033));
inv add_76_69_g1239 (.a(add_76_69_n_1038), .y(add_76_69_n_1037));
inv add_76_69_g1240 (.a(add_76_69_n_1039), .y(add_76_69_n_1040));
inv add_76_69_g1241 (.a(add_76_69_n_1042), .y(add_76_69_n_1041));
nand2 add_76_69_g1242 (.a(n_965), .b(v1_5_), .y(add_76_69_n_1044));
nand2 add_76_69_g1243 (.a(n_951), .b(v1_19_), .y(add_76_69_n_1046));
nand2 add_76_69_g1244 (.a(n_947), .b(v1_23_), .y(add_76_69_n_1047));
nor2 add_76_69_g1245 (.a(v1_6_), .b(v1_1_), .y(add_76_69_n_1001));
nand2 add_76_69_g1246 (.a(n_959), .b(v1_11_), .y(add_76_69_n_1003));
nand2 add_76_69_g1247 (.a(v1_27_), .b(v1_23_), .y(add_76_69_n_1048));
nand2 add_76_69_g1248 (.a(v1_8_), .b(v1_3_), .y(add_76_69_n_1051));
nand2 add_76_69_g1249 (.a(n_961), .b(v1_9_), .y(add_76_69_n_1007));
nand2 add_76_69_g1250 (.a(n_945), .b(v1_25_), .y(add_76_69_n_1009));
nand2 add_76_69_g1251 (.a(v1_6_), .b(v1_1_), .y(add_76_69_n_1010));
nand2 add_76_69_g1252 (.a(v1_29_), .b(v1_25_), .y(add_76_69_n_1012));
nand2 add_76_69_g1253 (.a(v1_5_), .b(v1_0_), .y(add_76_69_n_1013));
nor2 add_76_69_g1254 (.a(v1_7_), .b(v1_2_), .y(add_76_69_n_1015));
nand2 add_76_69_g1255 (.a(n_958), .b(v1_12_), .y(add_76_69_n_1017));
nand2 add_76_69_g1256 (.a(n_948), .b(v1_22_), .y(add_76_69_n_1018));
nor2 add_76_69_g1257 (.a(n_949), .b(v1_21_), .y(add_76_69_n_1019));
nand2 add_76_69_g1258 (.a(n_966), .b(v1_4_), .y(add_76_69_n_1021));
nor2 add_76_69_g1259 (.a(n_966), .b(v1_4_), .y(add_76_69_n_1023));
nand2 add_76_69_g1260 (.a(n_952), .b(v1_18_), .y(add_76_69_n_1025));
nor2 add_76_69_g1261 (.a(n_951), .b(v1_19_), .y(add_76_69_n_1026));
nand2 add_76_69_g1262 (.a(n_946), .b(v1_24_), .y(add_76_69_n_1060));
nor2 add_76_69_g1263 (.a(n_957), .b(v1_13_), .y(add_76_69_n_1028));
nor2 add_76_69_g1264 (.a(n_955), .b(v1_15_), .y(add_76_69_n_1030));
nand2 add_76_69_g1265 (.a(v1_7_), .b(v1_2_), .y(add_76_69_n_1032));
nor2 add_76_69_g1266 (.a(n_962), .b(v1_8_), .y(add_76_69_n_1034));
nand2 add_76_69_g1267 (.a(n_954), .b(v1_16_), .y(add_76_69_n_1036));
nor2 add_76_69_g1268 (.a(n_944), .b(v1_26_), .y(add_76_69_n_1038));
nor2 add_76_69_g1269 (.a(n_960), .b(v1_10_), .y(add_76_69_n_1039));
nor2 add_76_69_g1270 (.a(n_950), .b(v1_20_), .y(add_76_69_n_1042));
nor2 add_76_69_g1271 (.a(n_946), .b(v1_24_), .y(add_76_69_n_1043));
inv add_76_69_g1272 (.a(add_76_69_n_1110), .y(add_76_69_n_1066));
inv add_76_69_g1273 (.a(add_76_69_n_1111), .y(add_76_69_n_1067));
inv add_76_69_g1274 (.a(add_76_69_n_1114), .y(add_76_69_n_1068));
inv add_76_69_g1275 (.a(add_76_69_n_1070), .y(add_76_69_n_1069));
inv add_76_69_g1276 (.a(add_76_69_n_1117), .y(add_76_69_n_1071));
inv add_76_69_g1277 (.a(add_76_69_n_1119), .y(add_76_69_n_1072));
inv add_76_69_g1278 (.a(add_76_69_n_1075), .y(add_76_69_n_1076));
inv add_76_69_g1279 (.a(add_76_69_n_1081), .y(add_76_69_n_1080));
inv add_76_69_g1280 (.a(add_76_69_n_1083), .y(add_76_69_n_1082));
inv add_76_69_g1281 (.a(add_76_69_n_1087), .y(add_76_69_n_1086));
inv add_76_69_g1283 (.a(add_76_69_n_1093), .y(add_76_69_n_1092));
inv add_76_69_g1284 (.a(add_76_69_n_1095), .y(add_76_69_n_1094));
inv add_76_69_g1285 (.a(add_76_69_n_1098), .y(add_76_69_n_1097));
inv add_76_69_g1286 (.a(add_76_69_n_1100), .y(add_76_69_n_1099));
inv add_76_69_g1287 (.a(add_76_69_n_1103), .y(add_76_69_n_1102));
inv add_76_69_g1288 (.a(add_76_69_n_1107), .y(add_76_69_n_1106));
inv add_76_69_g1289 (.a(add_76_69_n_1108), .y(add_76_69_n_1109));
nand2 add_76_69_g1290 (.a(n_953), .b(v1_17_), .y(add_76_69_n_1110));
nand2 add_76_69_g1291 (.a(n_957), .b(v1_13_), .y(add_76_69_n_1111));
nand2 add_76_69_g1292 (.a(n_963), .b(v1_7_), .y(add_76_69_n_1114));
nand2 add_76_69_g1293 (.a(n_955), .b(v1_15_), .y(add_76_69_n_1070));
nand2 add_76_69_g1294 (.a(v1_30_), .b(v1_26_), .y(add_76_69_n_1117));
nand2 add_76_69_g1295 (.a(n_949), .b(v1_21_), .y(add_76_69_n_1119));
nor2 add_76_69_g1296 (.a(n_947), .b(v1_23_), .y(add_76_69_n_1073));
nor2 add_76_69_g1297 (.a(v1_8_), .b(v1_3_), .y(add_76_69_n_1074));
nor2 add_76_69_g1298 (.a(n_945), .b(v1_25_), .y(add_76_69_n_1075));
nor2 add_76_69_g1299 (.a(n_953), .b(v1_17_), .y(add_76_69_n_1077));
nor2 add_76_69_g1300 (.a(n_965), .b(v1_5_), .y(add_76_69_n_1078));
nor2 add_76_69_g1301 (.a(n_961), .b(v1_9_), .y(add_76_69_n_1079));
nand2 add_76_69_g1302 (.a(n_964), .b(v1_6_), .y(add_76_69_n_1081));
nor2 add_76_69_g1303 (.a(v1_29_), .b(v1_25_), .y(add_76_69_n_1083));
nor2 add_76_69_g1304 (.a(v1_30_), .b(v1_26_), .y(add_76_69_n_1084));
nand2 add_76_69_g1305 (.a(n_944), .b(v1_26_), .y(add_76_69_n_1085));
nor2 add_76_69_g1306 (.a(n_959), .b(v1_11_), .y(add_76_69_n_1087));
nand2 add_76_69_g1307 (.a(n_962), .b(v1_8_), .y(add_76_69_n_1088));
nor2 add_76_69_g1308 (.a(n_954), .b(v1_16_), .y(add_76_69_n_1090));
nor2 add_76_69_g1309 (.a(n_963), .b(v1_7_), .y(add_76_69_n_1091));
nand2 add_76_69_g1310 (.a(n_950), .b(v1_20_), .y(add_76_69_n_1093));
nand2 add_76_69_g1311 (.a(n_960), .b(v1_10_), .y(add_76_69_n_1095));
nor2 add_76_69_g1312 (.a(v1_27_), .b(v1_23_), .y(add_76_69_n_1096));
nand2 add_76_69_g1313 (.a(n_956), .b(v1_14_), .y(add_76_69_n_1098));
nand2 add_76_69_g1314 (.a(v1_28_), .b(v1_24_), .y(add_76_69_n_1100));
nor2 add_76_69_g1315 (.a(n_964), .b(v1_6_), .y(add_76_69_n_1101));
nor2 add_76_69_g1316 (.a(n_956), .b(v1_14_), .y(add_76_69_n_1103));
nor2 add_76_69_g1317 (.a(n_952), .b(v1_18_), .y(add_76_69_n_1104));
nor2 add_76_69_g1318 (.a(v1_28_), .b(v1_24_), .y(add_76_69_n_1105));
nor2 add_76_69_g1319 (.a(n_958), .b(v1_12_), .y(add_76_69_n_1107));
nor2 add_76_69_g1320 (.a(n_948), .b(v1_22_), .y(add_76_69_n_1108));
nand2 add_88_82_g1933 (.a(n_2993), .b(add_88_82_n_2235), .y(add_88_82_n_1889));
nand2 add_88_82_g1936 (.a(add_88_82_n_1896), .b(add_88_82_n_2145), .y(add_88_82_n_1893));
nand2 add_88_82_g1938 (.a(add_88_82_n_1900), .b(add_88_82_n_2283), .y(add_88_82_n_1896));
xor2 add_88_82_g1939 (.a(add_88_82_n_1905), .b(add_88_82_n_2126), .y(n_798));
nand2 add_88_82_g1941 (.a(add_88_82_n_1903), .b(add_88_82_n_2246), .y(add_88_82_n_1899));
nand2 add_88_82_g1942 (.a(add_88_82_n_1906), .b(add_88_82_n_2242), .y(add_88_82_n_1900));
xor2 add_88_82_g1943 (.a(add_88_82_n_1910), .b(add_88_82_n_2111), .y(n_825));
nand2 add_88_82_g1944 (.a(add_88_82_n_1910), .b(add_88_82_n_2170), .y(add_88_82_n_1903));
nand2 add_88_82_g1945 (.a(add_88_82_n_1911), .b(add_88_82_n_2155), .y(add_88_82_n_1905));
nand2 add_88_82_g1946 (.a(add_88_82_n_1913), .b(add_88_82_n_2287), .y(add_88_82_n_1906));
xor2 add_88_82_g1948 (.a(add_88_82_n_1921), .b(add_88_82_n_2127), .y(n_795));
nand2 add_88_82_g1950 (.a(add_88_82_n_1918), .b(add_88_82_n_2251), .y(add_88_82_n_1910));
nand2 add_88_82_g1951 (.a(add_88_82_n_1921), .b(add_88_82_n_2166), .y(add_88_82_n_1911));
nand2 add_88_82_g1952 (.a(add_88_82_n_1917), .b(add_88_82_n_2147), .y(add_88_82_n_1913));
nand2 add_88_82_g1955 (.a(add_88_82_n_1926), .b(add_88_82_n_2208), .y(add_88_82_n_1917));
nand2 add_88_82_g1956 (.a(add_88_82_n_1925), .b(add_88_82_n_2268), .y(add_88_82_n_1918));
nand2 add_88_82_g1957 (.a(add_88_82_n_1928), .b(add_88_82_n_2252), .y(add_88_82_n_1920));
nand2 add_88_82_g1958 (.a(add_88_82_n_1930), .b(add_88_82_n_2163), .y(add_88_82_n_1921));
nand2 add_88_82_g1962 (.a(add_88_82_n_1936), .b(add_88_82_n_2159), .y(add_88_82_n_1925));
nand2 add_88_82_g1963 (.a(add_88_82_n_1939), .b(add_88_82_n_2148), .y(add_88_82_n_1926));
nand2 add_88_82_g1964 (.a(add_88_82_n_1938), .b(add_88_82_n_2259), .y(add_88_82_n_1928));
nand2 add_88_82_g1965 (.a(add_88_82_n_1940), .b(add_88_82_n_2180), .y(add_88_82_n_1930));
nand2 add_88_82_g1966 (.a(add_88_82_n_1941), .b(add_88_82_n_2156), .y(add_88_82_n_1932));
xor2 add_88_82_g1968 (.a(add_88_82_n_1949), .b(add_88_82_n_2125), .y(n_801));
nand2 add_88_82_g1970 (.a(add_88_82_n_1945), .b(add_88_82_n_2164), .y(add_88_82_n_1936));
nand2 add_88_82_g1971 (.a(add_88_82_n_1947), .b(add_88_82_n_2161), .y(add_88_82_n_1938));
nand2 add_88_82_g1972 (.a(n_3975), .b(add_88_82_n_2005), .y(add_88_82_n_1939));
nand2 add_88_82_g1973 (.a(add_88_82_n_1950), .b(add_88_82_n_2253), .y(add_88_82_n_1940));
nand2 add_88_82_g1974 (.a(add_88_82_n_1952), .b(add_88_82_n_2172), .y(add_88_82_n_1941));
xor2 add_88_82_g1976 (.a(add_88_82_n_1960), .b(add_88_82_n_2129), .y(n_789));
nand2 add_88_82_g1977 (.a(n_3977), .b(add_88_82_n_2158), .y(add_88_82_n_1945));
nand2 add_88_82_g1979 (.a(add_88_82_n_1958), .b(add_88_82_n_2176), .y(add_88_82_n_1947));
nand2 add_88_82_g1980 (.a(add_88_82_n_1959), .b(add_88_82_n_2007), .y(add_88_82_n_1949));
nand2 add_88_82_g1981 (.a(add_88_82_n_1960), .b(add_88_82_n_2168), .y(add_88_82_n_1950));
nand2 add_88_82_g1982 (.a(add_88_82_n_1961), .b(add_88_82_n_2154), .y(add_88_82_n_1952));
xor2 add_88_82_g1984 (.a(add_88_82_n_1971), .b(add_88_82_n_2133), .y(n_777));
nand2 add_88_82_g1987 (.a(add_88_82_n_1965), .b(add_88_82_n_2247), .y(add_88_82_n_1958));
nand2 add_88_82_g1988 (.a(add_88_82_n_1968), .b(add_88_82_n_2035), .y(add_88_82_n_1959));
nand2 add_88_82_g1989 (.a(add_88_82_n_1969), .b(add_88_82_n_2249), .y(add_88_82_n_1960));
nand2 add_88_82_g1990 (.a(add_88_82_n_1971), .b(add_88_82_n_2178), .y(add_88_82_n_1961));
nand2 add_88_82_g1993 (.a(add_88_82_n_1973), .b(add_88_82_n_2263), .y(add_88_82_n_1965));
nand2 add_88_82_g1994 (.a(add_88_82_n_1977), .b(add_88_82_n_2004), .y(add_88_82_n_1967));
inv add_88_82_g1995 (.a(add_88_82_n_1969), .y(add_88_82_n_1968));
nand2 add_88_82_g1996 (.a(add_88_82_n_1974), .b(add_88_82_n_2174), .y(add_88_82_n_1969));
nand2 add_88_82_g1997 (.a(add_88_82_n_1975), .b(add_88_82_n_2245), .y(add_88_82_n_1971));
nand2 add_88_82_g1999 (.a(add_88_82_n_1982), .b(add_88_82_n_2257), .y(add_88_82_n_1973));
nand2 add_88_82_g2000 (.a(add_88_82_n_2372), .b(add_88_82_n_2003), .y(add_88_82_n_1974));
nand2 add_88_82_g2001 (.a(add_88_82_n_1981), .b(add_88_82_n_2265), .y(add_88_82_n_1975));
inv add_88_82_g2002 (.a(add_88_82_n_1978), .y(add_88_82_n_1977));
nor2 add_88_82_g2003 (.a(add_88_82_n_1982), .b(add_88_82_n_2045), .y(add_88_82_n_1978));
nand2 add_88_82_g2005 (.a(add_88_82_n_1985), .b(add_88_82_n_2244), .y(add_88_82_n_1981));
nor2 add_88_82_g2006 (.a(add_88_82_n_1987), .b(add_88_82_n_1993), .y(add_88_82_n_1982));
nand2 add_88_82_g2009 (.a(add_88_82_n_1989), .b(add_88_82_n_2254), .y(add_88_82_n_1985));
nor2 add_88_82_g2010 (.a(add_88_82_n_1988), .b(add_88_82_n_2011), .y(add_88_82_n_1987));
inv add_88_82_g2011 (.a(add_88_82_n_1989), .y(add_88_82_n_1988));
nand2 add_88_82_g2012 (.a(add_88_82_n_1991), .b(add_88_82_n_2293), .y(add_88_82_n_1989));
nand2 add_88_82_g2014 (.a(add_88_82_n_1994), .b(add_88_82_n_2238), .y(add_88_82_n_1991));
nor2 add_88_82_g2015 (.a(add_88_82_n_1996), .b(add_88_82_n_2152), .y(add_88_82_n_1993));
nand2 add_88_82_g2016 (.a(add_88_82_n_1997), .b(add_88_82_n_2271), .y(add_88_82_n_1994));
xor2 add_88_82_g2017 (.a(add_88_82_n_2001), .b(add_88_82_n_2131), .y(n_765));
nor2 add_88_82_g2018 (.a(add_88_82_n_1999), .b(add_88_82_n_2006), .y(add_88_82_n_1996));
nand2 add_88_82_g2019 (.a(add_88_82_n_2001), .b(add_88_82_n_2239), .y(add_88_82_n_1997));
nor2 add_88_82_g2020 (.a(add_88_82_n_2003), .b(add_88_82_n_2018), .y(add_88_82_n_1999));
nand2 add_88_82_g2021 (.a(add_88_82_n_2008), .b(add_88_82_n_2182), .y(add_88_82_n_2001));
nor2 add_88_82_g2023 (.a(add_88_82_n_2015), .b(add_88_82_n_2023), .y(add_88_82_n_2003));
nor2 add_88_82_g2024 (.a(add_88_82_n_2013), .b(add_88_82_n_2024), .y(add_88_82_n_2004));
nor2 add_88_82_g2025 (.a(add_88_82_n_2016), .b(add_88_82_n_2025), .y(add_88_82_n_2005));
inv add_88_82_g2026 (.a(add_88_82_n_2007), .y(add_88_82_n_2006));
nor2 add_88_82_g2027 (.a(add_88_82_n_2014), .b(add_88_82_n_2027), .y(add_88_82_n_2007));
nand2 add_88_82_g2028 (.a(add_88_82_n_2010), .b(add_88_82_n_2146), .y(add_88_82_n_2008));
nand2 add_88_82_g2029 (.a(n_2075), .b(add_88_82_n_2193), .y(add_88_82_n_2010));
nand2 add_88_82_g2030 (.a(add_88_82_n_2026), .b(add_88_82_n_2035), .y(add_88_82_n_2011));
nand2 add_88_82_g2031 (.a(add_88_82_n_2028), .b(add_88_82_n_2050), .y(add_88_82_n_2013));
nand2 add_88_82_g2032 (.a(add_88_82_n_2029), .b(add_88_82_n_2055), .y(add_88_82_n_2014));
nand2 add_88_82_g2033 (.a(add_88_82_n_2030), .b(add_88_82_n_2059), .y(add_88_82_n_2015));
nand2 add_88_82_g2034 (.a(add_88_82_n_2020), .b(add_88_82_n_2060), .y(add_88_82_n_2016));
nand2 add_88_82_g2036 (.a(add_88_82_n_2035), .b(add_88_82_n_2174), .y(add_88_82_n_2018));
nand2 add_88_82_g2037 (.a(add_88_82_n_2038), .b(add_88_82_n_2091), .y(add_88_82_n_2020));
nand2 add_88_82_g2039 (.a(add_88_82_n_2044), .b(add_88_82_n_2057), .y(add_88_82_n_2023));
nand2 add_88_82_g2040 (.a(add_88_82_n_2040), .b(add_88_82_n_2052), .y(add_88_82_n_2024));
nand2 add_88_82_g2041 (.a(add_88_82_n_2037), .b(add_88_82_n_2054), .y(add_88_82_n_2025));
nor2 add_88_82_g2042 (.a(add_88_82_n_2053), .b(add_88_82_n_2034), .y(add_88_82_n_2026));
nand2 add_88_82_g2043 (.a(add_88_82_n_2041), .b(add_88_82_n_2051), .y(add_88_82_n_2027));
nand2 add_88_82_g2044 (.a(add_88_82_n_2039), .b(add_88_82_n_2081), .y(add_88_82_n_2028));
nand2 add_88_82_g2045 (.a(add_88_82_n_2056), .b(add_88_82_n_2078), .y(add_88_82_n_2029));
nand2 add_88_82_g2046 (.a(add_88_82_n_2058), .b(add_88_82_n_2107), .y(add_88_82_n_2030));
inv add_88_82_g2050 (.a(add_88_82_n_2048), .y(add_88_82_n_2035));
nand2 add_88_82_g2051 (.a(add_88_82_n_2105), .b(add_88_82_n_2062), .y(add_88_82_n_2037));
nor2 add_88_82_g2052 (.a(add_88_82_n_2069), .b(add_88_82_n_2171), .y(add_88_82_n_2038));
nor2 add_88_82_g2053 (.a(add_88_82_n_2099), .b(add_88_82_n_2260), .y(add_88_82_n_2039));
nand2 add_88_82_g2054 (.a(add_88_82_n_2088), .b(add_88_82_n_2061), .y(add_88_82_n_2040));
nand2 add_88_82_g2055 (.a(add_88_82_n_2065), .b(add_88_82_n_2064), .y(add_88_82_n_2041));
nand2 add_88_82_g2056 (.a(add_88_82_n_2062), .b(add_88_82_n_2101), .y(add_88_82_n_2042));
nand2 add_88_82_g2057 (.a(add_88_82_n_2067), .b(add_88_82_n_2063), .y(add_88_82_n_2044));
nand2 add_88_82_g2058 (.a(add_88_82_n_2061), .b(add_88_82_n_2109), .y(add_88_82_n_2045));
nand2 add_88_82_g2059 (.a(add_88_82_n_2063), .b(add_88_82_n_2086), .y(add_88_82_n_2034));
nand2 add_88_82_g2060 (.a(add_88_82_n_2064), .b(add_88_82_n_2076), .y(add_88_82_n_2048));
nor2 add_88_82_g2062 (.a(add_88_82_n_2096), .b(add_88_82_n_2149), .y(add_88_82_n_2050));
nand2 add_88_82_g2063 (.a(add_88_82_n_2064), .b(add_88_82_n_2162), .y(add_88_82_n_2051));
nand2 add_88_82_g2064 (.a(add_88_82_n_2061), .b(add_88_82_n_2160), .y(add_88_82_n_2052));
nand2 add_88_82_g2065 (.a(add_88_82_n_2079), .b(add_88_82_n_2174), .y(add_88_82_n_2053));
nand2 add_88_82_g2066 (.a(add_88_82_n_2062), .b(add_88_82_n_2250), .y(add_88_82_n_2054));
nor2 add_88_82_g2067 (.a(add_88_82_n_2093), .b(add_88_82_n_2236), .y(add_88_82_n_2055));
nor2 add_88_82_g2068 (.a(add_88_82_n_2074), .b(add_88_82_n_2167), .y(add_88_82_n_2056));
nand2 add_88_82_g2069 (.a(add_88_82_n_2063), .b(add_88_82_n_2153), .y(add_88_82_n_2057));
nor2 add_88_82_g2070 (.a(add_88_82_n_2084), .b(add_88_82_n_2173), .y(add_88_82_n_2058));
nor2 add_88_82_g2071 (.a(add_88_82_n_2103), .b(add_88_82_n_2241), .y(add_88_82_n_2059));
nor2 add_88_82_g2072 (.a(add_88_82_n_2082), .b(add_88_82_n_2237), .y(add_88_82_n_2060));
nor2 add_88_82_g2073 (.a(add_88_82_n_2253), .b(add_88_82_n_2181), .y(add_88_82_n_2065));
nor2 add_88_82_g2074 (.a(add_88_82_n_2245), .b(add_88_82_n_2179), .y(add_88_82_n_2067));
nand2 add_88_82_g2075 (.a(add_88_82_n_2157), .b(add_88_82_n_2164), .y(add_88_82_n_2069));
nand2 add_88_82_g2078 (.a(add_88_82_n_2248), .b(add_88_82_n_2168), .y(add_88_82_n_2074));
nor2 add_88_82_g2079 (.a(add_88_82_n_2181), .b(add_88_82_n_2169), .y(add_88_82_n_2076));
nor2 add_88_82_g2080 (.a(add_88_82_n_2267), .b(add_88_82_n_2181), .y(add_88_82_n_2078));
nor2 add_88_82_g2081 (.a(add_88_82_n_2152), .b(add_88_82_n_2255), .y(add_88_82_n_2079));
nor2 add_88_82_g2082 (.a(add_88_82_n_2258), .b(add_88_82_n_2177), .y(add_88_82_n_2081));
nor2 add_88_82_g2083 (.a(add_88_82_n_2246), .b(add_88_82_n_2262), .y(add_88_82_n_2082));
nand2 add_88_82_g2084 (.a(add_88_82_n_2243), .b(add_88_82_n_2265), .y(add_88_82_n_2084));
nor2 add_88_82_g2085 (.a(add_88_82_n_2179), .b(add_88_82_n_2266), .y(add_88_82_n_2086));
nor2 add_88_82_g2086 (.a(add_88_82_n_2247), .b(add_88_82_n_2177), .y(add_88_82_n_2088));
nor2 add_88_82_g2087 (.a(add_88_82_n_2262), .b(add_88_82_n_2269), .y(add_88_82_n_2091));
nor2 add_88_82_g2088 (.a(add_88_82_n_2155), .b(add_88_82_n_2267), .y(add_88_82_n_2093));
nor2 add_88_82_g2089 (.a(add_88_82_n_2252), .b(add_88_82_n_2258), .y(add_88_82_n_2096));
nand2 add_88_82_g2090 (.a(add_88_82_n_2256), .b(add_88_82_n_2263), .y(add_88_82_n_2099));
nor2 add_88_82_g2091 (.a(add_88_82_n_2269), .b(add_88_82_n_2165), .y(add_88_82_n_2101));
nor2 add_88_82_g2092 (.a(add_88_82_n_2156), .b(add_88_82_n_2261), .y(add_88_82_n_2103));
nor2 add_88_82_g2093 (.a(add_88_82_n_2159), .b(add_88_82_n_2269), .y(add_88_82_n_2105));
nor2 add_88_82_g2094 (.a(add_88_82_n_2261), .b(add_88_82_n_2179), .y(add_88_82_n_2107));
nor2 add_88_82_g2095 (.a(add_88_82_n_2177), .b(add_88_82_n_2264), .y(add_88_82_n_2109));
xor2 add_88_82_g2096 (.a(n_681), .b(n_1286), .y(add_88_82_n_2110));
xor2 add_88_82_g2097 (.a(n_680), .b(n_1287), .y(add_88_82_n_2111));
nor2 add_88_82_g2098 (.a(add_88_82_n_2258), .b(add_88_82_n_2260), .y(add_88_82_n_2061));
nor2 add_88_82_g2099 (.a(add_88_82_n_2262), .b(add_88_82_n_2171), .y(add_88_82_n_2062));
nor2 add_88_82_g2100 (.a(add_88_82_n_2261), .b(add_88_82_n_2173), .y(add_88_82_n_2063));
nor2 add_88_82_g2101 (.a(add_88_82_n_2267), .b(add_88_82_n_2167), .y(add_88_82_n_2064));
xor2 add_88_82_g2102 (.a(n_666), .b(n_1301), .y(add_88_82_n_2116));
xor2 add_88_82_g2103 (.a(n_678), .b(n_1289), .y(add_88_82_n_2117));
xor2 add_88_82_g2104 (.a(n_677), .b(n_1290), .y(add_88_82_n_2118));
xor2 add_88_82_g2106 (.a(n_667), .b(n_3838), .y(add_88_82_n_2120));
xor2 add_88_82_g2107 (.a(n_676), .b(n_1291), .y(add_88_82_n_2121));
xor2 add_88_82_g2108 (.a(n_675), .b(n_1292), .y(add_88_82_n_2122));
xor2 add_88_82_g2109 (.a(n_674), .b(n_1293), .y(add_88_82_n_2123));
xor2 add_88_82_g2110 (.a(n_673), .b(n_1294), .y(add_88_82_n_2124));
xor2 add_88_82_g2111 (.a(n_672), .b(n_1295), .y(add_88_82_n_2125));
xor2 add_88_82_g2112 (.a(n_671), .b(n_1296), .y(add_88_82_n_2126));
xor2 add_88_82_g2113 (.a(n_670), .b(n_1297), .y(add_88_82_n_2127));
xor2 add_88_82_g2114 (.a(n_669), .b(n_1298), .y(add_88_82_n_2128));
xor2 add_88_82_g2115 (.a(n_668), .b(n_3814), .y(add_88_82_n_2129));
xor2 add_88_82_g2116 (.a(n_679), .b(n_1288), .y(add_88_82_n_2130));
xor2 add_88_82_g2117 (.a(n_660), .b(n_1307), .y(add_88_82_n_2131));
xor2 add_88_82_g2118 (.a(n_665), .b(n_1302), .y(add_88_82_n_2132));
xor2 add_88_82_g2119 (.a(n_664), .b(n_1303), .y(add_88_82_n_2133));
xor2 add_88_82_g2120 (.a(n_663), .b(n_1304), .y(add_88_82_n_2134));
xor2 add_88_82_g2121 (.a(n_662), .b(n_1305), .y(add_88_82_n_2135));
xor2 add_88_82_g2122 (.a(n_661), .b(n_1306), .y(add_88_82_n_2136));
xor2 add_88_82_g2123 (.a(n_659), .b(n_1308), .y(add_88_82_n_2137));
xor2 add_88_82_g2124 (.a(n_2080), .b(n_2070), .y(add_88_82_n_2138));
xor2 add_88_82_g2125 (.a(n_2065), .b(n_2066), .y(add_88_82_n_2139));
xor2 add_88_82_g2127 (.a(n_685), .b(n_1282), .y(add_88_82_n_2141));
xor2 add_88_82_g2128 (.a(n_684), .b(n_1283), .y(add_88_82_n_2142));
xor2 add_88_82_g2129 (.a(n_683), .b(n_1284), .y(add_88_82_n_2143));
xor2 add_88_82_g2130 (.a(n_682), .b(n_1285), .y(add_88_82_n_2144));
inv add_88_82_g2131 (.a(add_88_82_n_2185), .y(add_88_82_n_2145));
inv add_88_82_g2132 (.a(add_88_82_n_2189), .y(add_88_82_n_2146));
inv add_88_82_g2133 (.a(add_88_82_n_2190), .y(add_88_82_n_2147));
inv add_88_82_g2134 (.a(add_88_82_n_2199), .y(add_88_82_n_2148));
inv add_88_82_g2135 (.a(add_88_82_n_2202), .y(add_88_82_n_2149));
inv add_88_82_g2138 (.a(add_88_82_n_2154), .y(add_88_82_n_2153));
inv add_88_82_g2139 (.a(add_88_82_n_2158), .y(add_88_82_n_2157));
inv add_88_82_g2140 (.a(add_88_82_n_2161), .y(add_88_82_n_2160));
inv add_88_82_g2141 (.a(add_88_82_n_2163), .y(add_88_82_n_2162));
inv add_88_82_g2142 (.a(add_88_82_n_2165), .y(add_88_82_n_2164));
inv add_88_82_g2143 (.a(add_88_82_n_2167), .y(add_88_82_n_2166));
inv add_88_82_g2144 (.a(add_88_82_n_2169), .y(add_88_82_n_2168));
inv add_88_82_g2145 (.a(add_88_82_n_2171), .y(add_88_82_n_2170));
inv add_88_82_g2146 (.a(add_88_82_n_2173), .y(add_88_82_n_2172));
inv add_88_82_g2147 (.a(add_88_82_n_2231), .y(add_88_82_n_2174));
inv add_88_82_g2149 (.a(add_88_82_n_2177), .y(add_88_82_n_2176));
inv add_88_82_g2150 (.a(add_88_82_n_2179), .y(add_88_82_n_2178));
inv add_88_82_g2151 (.a(add_88_82_n_2181), .y(add_88_82_n_2180));
nand2 add_88_82_g2152 (.a(n_659), .b(n_1308), .y(add_88_82_n_2182));
nor2 add_88_82_g2153 (.a(n_685), .b(n_1282), .y(add_88_82_n_2185));
nand2 add_88_82_g2154 (.a(n_685), .b(n_1282), .y(add_88_82_n_2188));
nor2 add_88_82_g2155 (.a(n_659), .b(n_1308), .y(add_88_82_n_2189));
nor2 add_88_82_g2156 (.a(n_683), .b(n_1284), .y(add_88_82_n_2190));
nand2 add_88_82_g2157 (.a(n_2080), .b(n_2070), .y(add_88_82_n_2193));
nand2 add_88_82_g2158 (.a(n_686), .b(n_1281), .y(add_88_82_n_2196));
nor2 add_88_82_g2159 (.a(n_682), .b(n_1285), .y(add_88_82_n_2199));
nand2 add_88_82_g2160 (.a(n_676), .b(n_1291), .y(add_88_82_n_2202));
nand2 add_88_82_g2162 (.a(n_682), .b(n_1285), .y(add_88_82_n_2208));
nor2 add_88_82_g2165 (.a(n_672), .b(n_1295), .y(add_88_82_n_2152));
nand2 add_88_82_g2166 (.a(n_664), .b(n_1303), .y(add_88_82_n_2154));
nand2 add_88_82_g2167 (.a(n_670), .b(n_1297), .y(add_88_82_n_2155));
nand2 add_88_82_g2168 (.a(n_665), .b(n_1302), .y(add_88_82_n_2156));
nand2 add_88_82_g2169 (.a(n_677), .b(n_1290), .y(add_88_82_n_2158));
nand2 add_88_82_g2170 (.a(n_678), .b(n_1289), .y(add_88_82_n_2159));
nand2 add_88_82_g2171 (.a(n_674), .b(n_1293), .y(add_88_82_n_2161));
nand2 add_88_82_g2172 (.a(n_669), .b(n_1298), .y(add_88_82_n_2163));
nor2 add_88_82_g2173 (.a(n_678), .b(n_1289), .y(add_88_82_n_2165));
nor2 add_88_82_g2174 (.a(n_670), .b(n_1297), .y(add_88_82_n_2167));
nor2 add_88_82_g2175 (.a(n_668), .b(n_3814), .y(add_88_82_n_2169));
nor2 add_88_82_g2176 (.a(n_680), .b(n_1287), .y(add_88_82_n_2171));
nor2 add_88_82_g2177 (.a(n_665), .b(n_1302), .y(add_88_82_n_2173));
nor2 add_88_82_g2178 (.a(n_667), .b(n_3838), .y(add_88_82_n_2231));
nor2 add_88_82_g2180 (.a(n_674), .b(n_1293), .y(add_88_82_n_2177));
nor2 add_88_82_g2181 (.a(n_664), .b(n_1303), .y(add_88_82_n_2179));
nor2 add_88_82_g2182 (.a(n_669), .b(n_1298), .y(add_88_82_n_2181));
inv add_88_82_g2183 (.a(add_88_82_n_2270), .y(add_88_82_n_2235));
inv add_88_82_g2184 (.a(add_88_82_n_2274), .y(add_88_82_n_2236));
inv add_88_82_g2185 (.a(add_88_82_n_2277), .y(add_88_82_n_2237));
inv add_88_82_g2186 (.a(add_88_82_n_2280), .y(add_88_82_n_2238));
inv add_88_82_g2187 (.a(add_88_82_n_2286), .y(add_88_82_n_2239));
inv add_88_82_g2189 (.a(add_88_82_n_2289), .y(add_88_82_n_2241));
inv add_88_82_g2190 (.a(add_88_82_n_2292), .y(add_88_82_n_2242));
inv add_88_82_g2191 (.a(add_88_82_n_2244), .y(add_88_82_n_2243));
inv add_88_82_g2192 (.a(add_88_82_n_2249), .y(add_88_82_n_2248));
inv add_88_82_g2193 (.a(add_88_82_n_2251), .y(add_88_82_n_2250));
inv add_88_82_g2194 (.a(add_88_82_n_2255), .y(add_88_82_n_2254));
inv add_88_82_g2195 (.a(add_88_82_n_2257), .y(add_88_82_n_2256));
inv add_88_82_g2196 (.a(add_88_82_n_2260), .y(add_88_82_n_2259));
inv add_88_82_g2197 (.a(add_88_82_n_2264), .y(add_88_82_n_2263));
inv add_88_82_g2198 (.a(add_88_82_n_2266), .y(add_88_82_n_2265));
inv add_88_82_g2199 (.a(add_88_82_n_2269), .y(add_88_82_n_2268));
nor2 add_88_82_g2200 (.a(n_686), .b(n_1281), .y(add_88_82_n_2270));
nand2 add_88_82_g2201 (.a(n_660), .b(n_1307), .y(add_88_82_n_2271));
nand2 add_88_82_g2202 (.a(n_671), .b(n_1296), .y(add_88_82_n_2274));
nand2 add_88_82_g2203 (.a(n_681), .b(n_1286), .y(add_88_82_n_2277));
nor2 add_88_82_g2204 (.a(n_661), .b(n_1306), .y(add_88_82_n_2280));
nand2 add_88_82_g2205 (.a(n_684), .b(n_1283), .y(add_88_82_n_2283));
nor2 add_88_82_g2206 (.a(n_660), .b(n_1307), .y(add_88_82_n_2286));
nand2 add_88_82_g2207 (.a(n_683), .b(n_1284), .y(add_88_82_n_2287));
nor2 add_88_82_g2208 (.a(n_677), .b(n_1290), .y(add_88_82_n_2288));
nand2 add_88_82_g2209 (.a(n_666), .b(n_1301), .y(add_88_82_n_2289));
nor2 add_88_82_g2210 (.a(n_684), .b(n_1283), .y(add_88_82_n_2292));
nand2 add_88_82_g2211 (.a(n_661), .b(n_1306), .y(add_88_82_n_2293));
nand2 add_88_82_g2213 (.a(n_662), .b(n_1305), .y(add_88_82_n_2244));
nand2 add_88_82_g2214 (.a(n_663), .b(n_1304), .y(add_88_82_n_2245));
nand2 add_88_82_g2215 (.a(n_680), .b(n_1287), .y(add_88_82_n_2246));
nand2 add_88_82_g2216 (.a(n_673), .b(n_1294), .y(add_88_82_n_2247));
nand2 add_88_82_g2217 (.a(n_667), .b(n_3838), .y(add_88_82_n_2249));
nand2 add_88_82_g2218 (.a(n_679), .b(n_1288), .y(add_88_82_n_2251));
nand2 add_88_82_g2219 (.a(n_675), .b(n_1292), .y(add_88_82_n_2252));
nand2 add_88_82_g2220 (.a(n_668), .b(n_3814), .y(add_88_82_n_2253));
nor2 add_88_82_g2221 (.a(n_662), .b(n_1305), .y(add_88_82_n_2255));
nand2 add_88_82_g2222 (.a(n_672), .b(n_1295), .y(add_88_82_n_2257));
nor2 add_88_82_g2223 (.a(n_676), .b(n_1291), .y(add_88_82_n_2258));
nor2 add_88_82_g2224 (.a(n_675), .b(n_1292), .y(add_88_82_n_2260));
nor2 add_88_82_g2225 (.a(n_666), .b(n_1301), .y(add_88_82_n_2261));
nor2 add_88_82_g2226 (.a(n_681), .b(n_1286), .y(add_88_82_n_2262));
nor2 add_88_82_g2227 (.a(n_673), .b(n_1294), .y(add_88_82_n_2264));
nor2 add_88_82_g2228 (.a(n_663), .b(n_1304), .y(add_88_82_n_2266));
nor2 add_88_82_g2229 (.a(n_671), .b(n_1296), .y(add_88_82_n_2267));
nor2 add_88_82_g2230 (.a(n_679), .b(n_1288), .y(add_88_82_n_2269));
inv add_88_82_g2231 (.a(add_88_82_n_2371), .y(add_88_82_n_2372));
nor2 add_88_82_g2232 (.a(add_88_82_n_1985), .b(add_88_82_n_2034), .y(add_88_82_n_2371));
xor2 inc_add_77_23_g508 (.a(inc_add_77_23_n_412), .b(sum_31_), .y(n_1280));
xor2 inc_add_77_23_g509 (.a(inc_add_77_23_n_411), .b(sum_29_), .y(n_1282));
xor2 inc_add_77_23_g510 (.a(inc_add_77_23_n_413), .b(sum_23_), .y(n_1288));
xor2 inc_add_77_23_g511 (.a(inc_add_77_23_n_428), .b(inc_add_77_23_n_562), .y(n_1294));
xor2 inc_add_77_23_g512 (.a(inc_add_77_23_n_424), .b(inc_add_77_23_n_569), .y(n_1285));
xor2 inc_add_77_23_g513 (.a(inc_add_77_23_n_421), .b(inc_add_77_23_n_591), .y(n_1291));
xor2 inc_add_77_23_g514 (.a(inc_add_77_23_n_430), .b(sum_30_), .y(n_1281));
xor2 inc_add_77_23_g515 (.a(inc_add_77_23_n_431), .b(sum_27_), .y(n_1284));
xor2 inc_add_77_23_g516 (.a(inc_add_77_23_n_439), .b(sum_22_), .y(n_1289));
xor2 inc_add_77_23_g517 (.a(inc_add_77_23_n_440), .b(sum_19_), .y(n_1292));
xor2 inc_add_77_23_g518 (.a(inc_add_77_23_n_433), .b(sum_24_), .y(n_1287));
xor2 inc_add_77_23_g519 (.a(inc_add_77_23_n_426), .b(sum_28_), .y(n_1283));
xor2 inc_add_77_23_g520 (.a(inc_add_77_23_n_441), .b(sum_25_), .y(n_1286));
xor2 inc_add_77_23_g521 (.a(inc_add_77_23_n_422), .b(sum_21_), .y(n_1290));
xor2 inc_add_77_23_g522 (.a(inc_add_77_23_n_427), .b(sum_18_), .y(n_1293));
xor2 inc_add_77_23_g523 (.a(inc_add_77_23_n_453), .b(sum_9_), .y(n_1302));
xor2 inc_add_77_23_g524 (.a(inc_add_77_23_n_462), .b(sum_14_), .y(n_1297));
nor2 inc_add_77_23_g525 (.a(inc_add_77_23_n_432), .b(inc_add_77_23_n_470), .y(inc_add_77_23_n_411));
nor2 inc_add_77_23_g526 (.a(inc_add_77_23_n_435), .b(inc_add_77_23_n_445), .y(inc_add_77_23_n_412));
nor2 inc_add_77_23_g527 (.a(inc_add_77_23_n_421), .b(inc_add_77_23_n_512), .y(inc_add_77_23_n_413));
xor2 inc_add_77_23_g529 (.a(inc_add_77_23_n_444), .b(sum_16_), .y(n_1295));
xor2 inc_add_77_23_g531 (.a(inc_add_77_23_n_460), .b(sum_15_), .y(n_1296));
xor2 inc_add_77_23_g532 (.a(inc_add_77_23_n_454), .b(sum_13_), .y(n_1298));
xor2 inc_add_77_23_g533 (.a(inc_add_77_23_n_451), .b(sum_10_), .y(n_1301));
nor2 inc_add_77_23_g534 (.a(inc_add_77_23_n_445), .b(inc_add_77_23_n_476), .y(inc_add_77_23_n_422));
nand2 inc_add_77_23_g535 (.a(inc_add_77_23_n_446), .b(inc_add_77_23_n_444), .y(inc_add_77_23_n_424));
nor2 inc_add_77_23_g536 (.a(inc_add_77_23_n_443), .b(inc_add_77_23_n_445), .y(inc_add_77_23_n_426));
nor2 inc_add_77_23_g537 (.a(inc_add_77_23_n_445), .b(inc_add_77_23_n_524), .y(inc_add_77_23_n_427));
nand2 inc_add_77_23_g538 (.a(inc_add_77_23_n_444), .b(sum_16_), .y(inc_add_77_23_n_428));
nor2 inc_add_77_23_g539 (.a(inc_add_77_23_n_458), .b(inc_add_77_23_n_445), .y(inc_add_77_23_n_430));
nor2 inc_add_77_23_g540 (.a(inc_add_77_23_n_455), .b(inc_add_77_23_n_445), .y(inc_add_77_23_n_431));
nand2 inc_add_77_23_g541 (.a(inc_add_77_23_n_444), .b(inc_add_77_23_n_491), .y(inc_add_77_23_n_421));
inv inc_add_77_23_g542 (.a(inc_add_77_23_n_433), .y(inc_add_77_23_n_432));
xor2 inc_add_77_23_g543 (.a(inc_add_77_23_n_486), .b(sum_6_), .y(n_1305));
nand2 inc_add_77_23_g544 (.a(inc_add_77_23_n_442), .b(inc_add_77_23_n_506), .y(inc_add_77_23_n_435));
mux2 inc_add_77_23_g545 (.a(n_3804), .b(inc_add_77_23_n_465), .sel(sum_8_), .y(n_1303));
xor2 inc_add_77_23_g546 (.a(inc_add_77_23_n_487), .b(sum_7_), .y(n_1304));
xor2 inc_add_77_23_g547 (.a(inc_add_77_23_n_478), .b(inc_add_77_23_n_585), .y(n_1306));
nor2 inc_add_77_23_g548 (.a(inc_add_77_23_n_445), .b(inc_add_77_23_n_484), .y(inc_add_77_23_n_439));
nor2 inc_add_77_23_g549 (.a(inc_add_77_23_n_445), .b(inc_add_77_23_n_517), .y(inc_add_77_23_n_440));
nor2 inc_add_77_23_g550 (.a(inc_add_77_23_n_448), .b(inc_add_77_23_n_445), .y(inc_add_77_23_n_441));
nor2 inc_add_77_23_g551 (.a(inc_add_77_23_n_445), .b(inc_add_77_23_n_463), .y(inc_add_77_23_n_433));
inv inc_add_77_23_g552 (.a(inc_add_77_23_n_443), .y(inc_add_77_23_n_442));
inv inc_add_77_23_g553 (.a(inc_add_77_23_n_444), .y(inc_add_77_23_n_445));
nor2 inc_add_77_23_g554 (.a(inc_add_77_23_n_463), .b(inc_add_77_23_n_544), .y(inc_add_77_23_n_446));
nand2 inc_add_77_23_g555 (.a(inc_add_77_23_n_464), .b(sum_24_), .y(inc_add_77_23_n_448));
nand2 inc_add_77_23_g556 (.a(inc_add_77_23_n_464), .b(inc_add_77_23_n_490), .y(inc_add_77_23_n_443));
nor2 inc_add_77_23_g557 (.a(n_3804), .b(inc_add_77_23_n_526), .y(inc_add_77_23_n_451));
nor2 inc_add_77_23_g558 (.a(n_3804), .b(inc_add_77_23_n_593), .y(inc_add_77_23_n_453));
nor2 inc_add_77_23_g559 (.a(n_4135), .b(n_3804), .y(inc_add_77_23_n_454));
nor2 inc_add_77_23_g560 (.a(inc_add_77_23_n_469), .b(n_3804), .y(inc_add_77_23_n_444));
nand2 inc_add_77_23_g561 (.a(inc_add_77_23_n_464), .b(inc_add_77_23_n_498), .y(inc_add_77_23_n_455));
xor2 inc_add_77_23_g562 (.a(inc_add_77_23_n_494), .b(sum_4_), .y(n_1307));
xor2 inc_add_77_23_g563 (.a(inc_add_77_23_n_520), .b(sum_3_), .y(n_1308));
nand2 inc_add_77_23_g564 (.a(inc_add_77_23_n_483), .b(inc_add_77_23_n_464), .y(inc_add_77_23_n_458));
nor2 inc_add_77_23_g566 (.a(inc_add_77_23_n_485), .b(n_3804), .y(inc_add_77_23_n_460));
nor2 inc_add_77_23_g568 (.a(inc_add_77_23_n_482), .b(n_3804), .y(inc_add_77_23_n_462));
inv inc_add_77_23_g569 (.a(inc_add_77_23_n_463), .y(inc_add_77_23_n_464));
inv inc_add_77_23_g570 (.a(n_3804), .y(inc_add_77_23_n_465));
nand2 inc_add_77_23_g571 (.a(inc_add_77_23_n_502), .b(inc_add_77_23_n_492), .y(inc_add_77_23_n_469));
nand2 inc_add_77_23_g572 (.a(inc_add_77_23_n_490), .b(sum_28_), .y(inc_add_77_23_n_470));
nand2 inc_add_77_23_g574 (.a(inc_add_77_23_n_491), .b(sum_20_), .y(inc_add_77_23_n_476));
nand2 inc_add_77_23_g575 (.a(inc_add_77_23_n_494), .b(sum_4_), .y(inc_add_77_23_n_478));
nand2 inc_add_77_23_g576 (.a(inc_add_77_23_n_501), .b(inc_add_77_23_n_491), .y(inc_add_77_23_n_463));
nand2 inc_add_77_23_g579 (.a(inc_add_77_23_n_492), .b(inc_add_77_23_n_545), .y(inc_add_77_23_n_482));
nor2 inc_add_77_23_g580 (.a(inc_add_77_23_n_489), .b(inc_add_77_23_n_522), .y(inc_add_77_23_n_483));
nand2 inc_add_77_23_g581 (.a(inc_add_77_23_n_491), .b(inc_add_77_23_n_540), .y(inc_add_77_23_n_484));
nand2 inc_add_77_23_g582 (.a(inc_add_77_23_n_515), .b(inc_add_77_23_n_492), .y(inc_add_77_23_n_485));
nor2 inc_add_77_23_g583 (.a(inc_add_77_23_n_495), .b(inc_add_77_23_n_543), .y(inc_add_77_23_n_486));
nor2 inc_add_77_23_g584 (.a(inc_add_77_23_n_510), .b(inc_add_77_23_n_495), .y(inc_add_77_23_n_487));
inv inc_add_77_23_g585 (.a(inc_add_77_23_n_490), .y(inc_add_77_23_n_489));
inv inc_add_77_23_g586 (.a(inc_add_77_23_n_492), .y(inc_add_77_23_n_493));
inv inc_add_77_23_g587 (.a(inc_add_77_23_n_494), .y(inc_add_77_23_n_495));
nor2 inc_add_77_23_g588 (.a(inc_add_77_23_n_530), .b(inc_add_77_23_n_543), .y(inc_add_77_23_n_496));
nor2 inc_add_77_23_g589 (.a(inc_add_77_23_n_544), .b(inc_add_77_23_n_569), .y(inc_add_77_23_n_498));
nor2 inc_add_77_23_g590 (.a(inc_add_77_23_n_528), .b(inc_add_77_23_n_541), .y(inc_add_77_23_n_501));
nor2 inc_add_77_23_g591 (.a(inc_add_77_23_n_532), .b(inc_add_77_23_n_546), .y(inc_add_77_23_n_502));
nor2 inc_add_77_23_g592 (.a(inc_add_77_23_n_551), .b(inc_add_77_23_n_544), .y(inc_add_77_23_n_490));
nor2 inc_add_77_23_g593 (.a(inc_add_77_23_n_547), .b(inc_add_77_23_n_524), .y(inc_add_77_23_n_491));
nor2 inc_add_77_23_g594 (.a(inc_add_77_23_n_553), .b(inc_add_77_23_n_526), .y(inc_add_77_23_n_492));
nor2 inc_add_77_23_g595 (.a(inc_add_77_23_n_549), .b(inc_add_77_23_n_527), .y(inc_add_77_23_n_494));
nor2 inc_add_77_23_g596 (.a(inc_add_77_23_n_522), .b(inc_add_77_23_n_581), .y(inc_add_77_23_n_506));
nand2 inc_add_77_23_g597 (.a(inc_add_77_23_n_525), .b(sum_10_), .y(inc_add_77_23_n_508));
nand2 inc_add_77_23_g598 (.a(inc_add_77_23_n_542), .b(sum_6_), .y(inc_add_77_23_n_510));
nand2 inc_add_77_23_g599 (.a(inc_add_77_23_n_540), .b(sum_22_), .y(inc_add_77_23_n_512));
nor2 inc_add_77_23_g600 (.a(inc_add_77_23_n_546), .b(inc_add_77_23_n_572), .y(inc_add_77_23_n_515));
nand2 inc_add_77_23_g601 (.a(inc_add_77_23_n_523), .b(sum_18_), .y(inc_add_77_23_n_517));
nor2 inc_add_77_23_g603 (.a(inc_add_77_23_n_527), .b(inc_add_77_23_n_566), .y(inc_add_77_23_n_520));
inv inc_add_77_23_g604 (.a(inc_add_77_23_n_524), .y(inc_add_77_23_n_523));
inv inc_add_77_23_g605 (.a(inc_add_77_23_n_526), .y(inc_add_77_23_n_525));
nand2 inc_add_77_23_g606 (.a(sum_23_), .b(sum_22_), .y(inc_add_77_23_n_528));
nand2 inc_add_77_23_g607 (.a(sum_7_), .b(sum_6_), .y(inc_add_77_23_n_530));
nand2 inc_add_77_23_g608 (.a(sum_15_), .b(sum_14_), .y(inc_add_77_23_n_532));
nand2 inc_add_77_23_g609 (.a(sum_29_), .b(sum_28_), .y(inc_add_77_23_n_522));
nand2 inc_add_77_23_g610 (.a(sum_17_), .b(sum_16_), .y(inc_add_77_23_n_524));
nand2 inc_add_77_23_g611 (.a(sum_9_), .b(sum_8_), .y(inc_add_77_23_n_526));
nand2 inc_add_77_23_g612 (.a(sum_1_), .b(sum_0_), .y(inc_add_77_23_n_527));
inv inc_add_77_23_g613 (.a(inc_add_77_23_n_541), .y(inc_add_77_23_n_540));
inv inc_add_77_23_g614 (.a(inc_add_77_23_n_543), .y(inc_add_77_23_n_542));
inv inc_add_77_23_g615 (.a(inc_add_77_23_n_546), .y(inc_add_77_23_n_545));
nand2 inc_add_77_23_g616 (.a(sum_19_), .b(sum_18_), .y(inc_add_77_23_n_547));
nand2 inc_add_77_23_g617 (.a(sum_3_), .b(sum_2_), .y(inc_add_77_23_n_549));
nand2 inc_add_77_23_g618 (.a(sum_27_), .b(sum_26_), .y(inc_add_77_23_n_551));
nand2 inc_add_77_23_g619 (.a(sum_11_), .b(sum_10_), .y(inc_add_77_23_n_553));
nand2 inc_add_77_23_g620 (.a(sum_21_), .b(sum_20_), .y(inc_add_77_23_n_541));
nand2 inc_add_77_23_g621 (.a(sum_5_), .b(sum_4_), .y(inc_add_77_23_n_543));
nand2 inc_add_77_23_g622 (.a(sum_25_), .b(sum_24_), .y(inc_add_77_23_n_544));
nand2 inc_add_77_23_g623 (.a(sum_13_), .b(sum_12_), .y(inc_add_77_23_n_546));
inv inc_add_77_23_g624 (.a(sum_17_), .y(inc_add_77_23_n_562));
inv inc_add_77_23_g625 (.a(sum_2_), .y(inc_add_77_23_n_566));
inv inc_add_77_23_g626 (.a(sum_26_), .y(inc_add_77_23_n_569));
inv inc_add_77_23_g627 (.a(sum_14_), .y(inc_add_77_23_n_572));
inv inc_add_77_23_g628 (.a(sum_30_), .y(inc_add_77_23_n_581));
inv inc_add_77_23_g629 (.a(sum_5_), .y(inc_add_77_23_n_585));
inv inc_add_77_23_g630 (.a(sum_20_), .y(inc_add_77_23_n_591));
inv inc_add_77_23_g631 (.a(sum_8_), .y(inc_add_77_23_n_593));
nor2 g2 (.a(n_1312), .b(n_3891), .y(n_1313));
nand2 g6451 (.a(n_2853), .b(n_2846), .y(n_1312));
nand2 add_88_21_g6452 (.a(n_1314), .b(n_2853), .y(n_1315));
inv add_88_21_g6453 (.a(n_3891), .y(n_1314));
nor2 add_76_21_g6455 (.a(n_1557), .b(v0_21_), .y(n_1322));
nand2 add_76_21_g6461 (.a(n_1557), .b(v0_21_), .y(n_1323));
nand2 add_76_21_g6468 (.a(n_2564), .b(v0_19_), .y(n_1330));
xor2 add_88_69_g1538__6485 (.a(n_1345), .b(n_1346), .y(n_1347));
xor2 add_88_82_g6486 (.a(add_88_82_n_1939), .b(add_88_82_n_2144), .y(n_1345));
nand2 add_88_69_g1778__6487 (.a(add_88_69_n_1717), .b(add_88_69_n_1669), .y(n_1346));
nor2 add_88_69_g1545__6488 (.a(n_3597), .b(add_88_69_n_1262), .y(n_1348));
xor2 add_88_69_g1535__6499 (.a(n_1359), .b(n_1360), .y(n_1361));
xor2 add_88_82_g6500 (.a(add_88_82_n_1896), .b(add_88_82_n_2141), .y(n_1359));
nand2 add_88_69_g6501 (.a(add_88_69_n_1705), .b(add_88_69_n_1715), .y(n_1360));
nor2 add_88_69_g1561__6502 (.a(add_88_69_n_1298), .b(add_88_69_n_1265), .y(n_1362));
nand2 add_76_21_g6517 (.a(n_2875), .b(v0_5_), .y(n_1379));
nand2 add_76_21_g6524 (.a(n_2300), .b(v0_13_), .y(n_1386));
xor2 add_88_69_g1528__6527 (.a(n_1387), .b(n_1388), .y(n_1389));
xor2 add_88_82_g6528 (.a(add_88_82_n_1925), .b(add_88_82_n_2130), .y(n_1387));
nor2 add_88_69_g6529 (.a(add_88_69_n_1634), .b(n_2587), .y(n_1388));
nand2 add_88_21_g6531 (.a(n_3638), .b(v1_23_), .y(n_1393));
nand2 add_76_21_g6538 (.a(n_2278), .b(v0_15_), .y(n_1400));
nand2 add_76_21_g6545 (.a(n_2289), .b(v0_14_), .y(n_1407));
nand2 add_76_21_g6552 (.a(n_2341), .b(v0_12_), .y(n_1414));
nand2 add_76_21_g6559 (.a(n_2352), .b(v0_11_), .y(n_1421));
nand2 add_76_21_g6566 (.a(n_3688), .b(v0_10_), .y(n_1428));
nand2 add_76_21_g6580 (.a(n_2718), .b(v0_7_), .y(n_1442));
xor2 add_76_82_g6582 (.a(n_1445), .b(n_1446), .y(n_1447));
xor2 add_76_69_g6583 (.a(n_1443), .b(n_1444), .y(n_1445));
nor2 add_76_82_g6584 (.a(add_76_82_n_1194), .b(add_76_82_n_1277), .y(n_1443));
nor2 add_76_69_g6585 (.a(add_76_69_n_1067), .b(add_76_69_n_1028), .y(n_1444));
nand2 add_76_69_g6586 (.a(add_76_69_n_714), .b(add_76_69_n_690), .y(n_1446));
xor2 g6445__6588 (.a(n_1451), .b(n_1452), .y(n_1453));
xor2 add_88_69_g1526__6589 (.a(n_1449), .b(n_1450), .y(n_1451));
xor2 add_88_82_g6590 (.a(add_88_82_n_1899), .b(add_88_82_n_2110), .y(n_1449));
nor2 add_88_69_g6591 (.a(add_88_69_n_1699), .b(add_88_69_n_1647), .y(n_1450));
nand2 add_88_69_g1549__6592 (.a(add_88_69_n_1318), .b(add_88_69_n_1259), .y(n_1452));
nand2 add_88_69_g1542__6599 (.a(add_88_69_n_1290), .b(add_88_69_n_1274), .y(n_1459));
xor2 add_76_69_g6603 (.a(n_1463), .b(n_1464), .y(n_1465));
nand2 add_76_82_g6604 (.a(add_76_82_n_1269), .b(add_76_82_n_1225), .y(n_1463));
nand2 add_76_69_g6605 (.a(add_76_69_n_1070), .b(add_76_69_n_1029), .y(n_1464));
xor2 add_76_82_g6608 (.a(n_1471), .b(n_1472), .y(n_1473));
xor2 add_76_69_g6609 (.a(n_1469), .b(n_1470), .y(n_1471));
nand2 add_76_82_g6610 (.a(add_76_82_n_1279), .b(add_76_82_n_1229), .y(n_1469));
nand2 add_76_69_g6611 (.a(add_76_69_n_1098), .b(add_76_69_n_1102), .y(n_1470));
nor2 add_76_69_g6612 (.a(add_76_69_n_710), .b(add_76_69_n_697), .y(n_1472));
xor2 add_76_82_g6614 (.a(n_1477), .b(n_1478), .y(n_1479));
xor2 add_76_69_g6615 (.a(n_1475), .b(n_1476), .y(n_1477));
nand2 add_76_82_g6616 (.a(add_76_82_n_1206), .b(add_76_82_n_1235), .y(n_1475));
nand2 add_76_69_g6617 (.a(add_76_69_n_1017), .b(add_76_69_n_1106), .y(n_1476));
nor2 add_76_69_g6618 (.a(add_76_69_n_698), .b(add_76_69_n_745), .y(n_1478));
xor2 add_88_69_g1530__6621 (.a(n_1481), .b(n_3926), .y(n_1483));
xor2 add_88_82_g6622 (.a(add_88_82_n_1967), .b(add_88_82_n_2118), .y(n_1481));
nand2 add_88_69_g1544__6624 (.a(add_88_69_n_1268), .b(add_88_69_n_1327), .y(n_1484));
nand2 add_88_21_g6625 (.a(n_3300), .b(v1_21_), .y(n_1487));
xor2 add_76_69_g6628 (.a(n_1488), .b(n_1489), .y(n_1490));
nand2 add_76_82_g6629 (.a(add_76_82_n_1199), .b(add_76_82_n_1294), .y(n_1488));
nand2 add_76_69_g6630 (.a(add_76_69_n_1003), .b(add_76_69_n_1086), .y(n_1489));
xor2 add_76_82_g6633 (.a(n_1496), .b(n_1497), .y(n_1498));
xor2 add_76_69_g6634 (.a(n_1494), .b(n_1495), .y(n_1496));
nor2 add_76_82_g6635 (.a(add_76_82_n_1227), .b(add_76_82_n_1237), .y(n_1494));
nor2 add_76_69_g6636 (.a(add_76_69_n_1094), .b(add_76_69_n_1039), .y(n_1495));
nand2 add_76_69_g6637 (.a(add_76_69_n_692), .b(add_76_69_n_839), .y(n_1497));
xor2 add_76_82_g6639 (.a(n_1502), .b(n_1503), .y(n_1504));
xor2 add_76_69_g6640 (.a(n_1500), .b(n_1501), .y(n_1502));
nor2 add_76_82_g6641 (.a(add_76_82_n_1266), .b(add_76_82_n_1223), .y(n_1500));
nor2 add_76_69_g6642 (.a(add_76_69_n_1006), .b(add_76_69_n_1079), .y(n_1501));
nand2 add_76_69_g6643 (.a(add_76_69_n_683), .b(add_76_69_n_1088), .y(n_1503));
nand2 add_76_21_g6644 (.a(n_1510), .b(v0_6_), .y(n_1511));
xor2 g6423__6645 (.a(n_1508), .b(n_1509), .y(n_1510));
xor2 add_76_82_g6646 (.a(n_2941), .b(n_1507), .y(n_1508));
nor2 add_76_82_g6648 (.a(add_76_82_n_1289), .b(add_76_82_n_1231), .y(n_1507));
nand2 add_76_82_g6649 (.a(n_3911), .b(add_76_82_n_1059), .y(n_1509));
nor2 add_76_21_g6650 (.a(n_1510), .b(v0_6_), .y(n_1512));
xor2 add_76_82_g6652 (.a(n_1515), .b(n_1516), .y(n_1517));
xor2 add_76_69_g6653 (.a(n_1513), .b(n_1514), .y(n_1515));
nor2 add_76_82_g6654 (.a(add_76_82_n_1264), .b(add_76_82_n_1224), .y(n_1513));
nor2 add_76_69_g6655 (.a(add_76_69_n_1068), .b(add_76_69_n_1091), .y(n_1514));
nand2 add_76_69_g6656 (.a(add_76_69_n_771), .b(add_76_69_n_742), .y(n_1516));
xor2 add_76_69_g6666 (.a(n_1526), .b(n_1527), .y(n_1528));
nand2 add_76_82_g6667 (.a(add_76_82_n_1263), .b(add_76_82_n_1274), .y(n_1526));
nor2 add_76_69_g6668 (.a(add_76_69_n_1066), .b(add_76_69_n_1077), .y(n_1527));
xor2 add_88_69_g1536__6678 (.a(n_1538), .b(n_1539), .y(n_1540));
xor2 add_88_82_g6679 (.a(add_88_82_n_1938), .b(add_88_82_n_2122), .y(n_1538));
nor2 add_88_69_g6680 (.a(add_88_69_n_1631), .b(add_88_69_n_1650), .y(n_1539));
nand2 add_88_69_g1560__6681 (.a(add_88_69_n_1276), .b(add_88_69_n_1380), .y(n_1541));
nand2 add_88_21_g6682 (.a(n_3293), .b(v1_19_), .y(n_1544));
nand2 add_76_21_g6683 (.a(n_1631), .b(v0_20_), .y(n_1550));
nor2 add_76_82_g6688 (.a(add_76_82_n_847), .b(add_76_82_n_936), .y(n_1548));
nor2 add_76_21_g6689 (.a(n_1631), .b(v0_20_), .y(n_1551));
xor2 g6409__6690 (.a(n_1556), .b(n_2219), .y(n_1557));
xor2 add_76_82_g6691 (.a(n_1554), .b(n_1555), .y(n_1556));
xor2 add_76_69_g6692 (.a(n_1552), .b(n_1553), .y(n_1554));
nor2 add_76_82_g6693 (.a(add_76_82_n_1261), .b(add_76_82_n_1286), .y(n_1552));
nor2 add_76_69_g6694 (.a(add_76_69_n_1072), .b(add_76_69_n_1019), .y(n_1553));
nand2 add_76_69_g6695 (.a(add_76_69_n_654), .b(add_76_69_n_711), .y(n_1555));
nor2 add_76_21_g6696 (.a(n_1644), .b(v0_23_), .y(n_1563));
nand2 add_76_82_g6701 (.a(add_76_82_n_848), .b(add_76_82_n_910), .y(n_1561));
nand2 add_76_21_g6702 (.a(n_1644), .b(v0_23_), .y(n_1564));
xor2 add_76_69_g6712 (.a(n_1572), .b(n_1573), .y(n_1574));
nor2 add_76_82_g6713 (.a(add_76_82_n_1201), .b(add_76_82_n_1222), .y(n_1572));
nor2 add_76_69_g6714 (.a(add_76_69_n_998), .b(add_76_69_n_1026), .y(n_1573));
xor2 add_88_69_g1529__6718 (.a(n_1578), .b(n_1579), .y(n_1580));
xor2 add_88_82_g6719 (.a(add_88_82_n_1945), .b(add_88_82_n_2117), .y(n_1578));
nand2 add_88_69_g6720 (.a(n_3574), .b(n_2841), .y(n_1579));
nand2 add_88_21_g6722 (.a(n_3727), .b(v1_22_), .y(n_1584));
nand2 add_88_21_g6723 (.a(n_1589), .b(v1_20_), .y(n_1590));
xor2 g2621__6724 (.a(n_1587), .b(n_1588), .y(n_1589));
xor2 add_88_69_g1525__6725 (.a(n_1585), .b(n_1586), .y(n_1587));
xor2 add_88_82_g6726 (.a(add_88_82_n_1920), .b(add_88_82_n_2121), .y(n_1585));
nand2 add_88_69_g6727 (.a(n_2520), .b(add_88_69_n_1741), .y(n_1586));
nor2 add_88_69_g1550__6728 (.a(add_88_69_n_1272), .b(add_88_69_n_1366), .y(n_1588));
nor2 add_88_21_g6729 (.a(n_1589), .b(v1_20_), .y(n_1591));
nor2 add_88_21_g6730 (.a(n_1596), .b(v1_18_), .y(n_1597));
xor2 g6449__6731 (.a(n_1594), .b(n_1595), .y(n_1596));
xor2 add_88_69_g1533__6732 (.a(n_1592), .b(n_1593), .y(n_1594));
xor2 add_88_82_g6733 (.a(add_88_82_n_1958), .b(add_88_82_n_2123), .y(n_1592));
nor2 add_88_69_g6734 (.a(add_88_69_n_1659), .b(add_88_69_n_1740), .y(n_1593));
nand2 add_88_69_g1540__6735 (.a(add_88_69_n_1261), .b(n_3887), .y(n_1595));
nand2 add_88_21_g6736 (.a(n_1596), .b(v1_18_), .y(n_1598));
nor2 add_76_21_g6743 (.a(n_1656), .b(v0_24_), .y(n_1605));
xor2 add_76_69_g6746 (.a(n_1606), .b(n_1607), .y(n_1608));
nor2 add_76_82_g6747 (.a(add_76_82_n_1260), .b(add_76_82_n_1284), .y(n_1606));
nor2 add_76_69_g6748 (.a(add_76_69_n_1008), .b(add_76_69_n_1075), .y(n_1607));
nor2 add_88_21_g6757 (.a(n_1623), .b(v1_17_), .y(n_1624));
xor2 g6389__6758 (.a(n_1621), .b(n_1622), .y(n_1623));
xor2 add_88_69_g1534__6759 (.a(n_1619), .b(n_1620), .y(n_1621));
xor2 add_88_82_g6760 (.a(add_88_82_n_1973), .b(add_88_82_n_2124), .y(n_1619));
nand2 add_88_69_g6761 (.a(add_88_69_n_1633), .b(add_88_69_n_1656), .y(n_1620));
nor2 add_88_69_g1546__6762 (.a(add_88_69_n_1328), .b(add_88_69_n_1263), .y(n_1622));
nand2 add_88_21_g6763 (.a(n_1623), .b(v1_17_), .y(n_1625));
xor2 g6410__6764 (.a(n_1630), .b(n_1548), .y(n_1631));
xor2 add_76_82_g6765 (.a(n_1628), .b(n_1629), .y(n_1630));
xor2 add_76_69_g6766 (.a(n_1626), .b(n_1627), .y(n_1628));
nand2 add_76_82_g6767 (.a(add_76_82_n_1217), .b(add_76_82_n_1297), .y(n_1626));
nand2 add_76_69_g6768 (.a(add_76_69_n_1093), .b(add_76_69_n_1041), .y(n_1627));
nor2 add_76_69_g6769 (.a(add_76_69_n_658), .b(add_76_69_n_743), .y(n_1629));
nor2 add_76_21_g6770 (.a(n_1636), .b(v0_22_), .y(n_1637));
xor2 g6408__6771 (.a(n_2230), .b(n_1635), .y(n_1636));
nand2 add_76_82_g6774 (.a(add_76_82_n_1215), .b(add_76_82_n_1301), .y(n_1633));
nor2 add_76_82_g6775 (.a(add_76_82_n_846), .b(add_76_82_n_904), .y(n_1635));
nand2 add_76_21_g6776 (.a(n_1636), .b(v0_22_), .y(n_1638));
xor2 g6407__6777 (.a(n_1643), .b(n_1561), .y(n_1644));
xor2 add_76_82_g6778 (.a(n_1641), .b(n_1642), .y(n_1643));
xor2 add_76_69_g6779 (.a(n_1639), .b(n_1640), .y(n_1641));
nor2 add_76_82_g6780 (.a(add_76_82_n_1200), .b(add_76_82_n_1204), .y(n_1639));
nor2 add_76_69_g6781 (.a(add_76_69_n_999), .b(add_76_69_n_1073), .y(n_1640));
nand2 add_76_69_g6782 (.a(add_76_69_n_659), .b(add_76_69_n_717), .y(n_1642));
xor2 add_76_69_g6785 (.a(n_1645), .b(n_1646), .y(n_1647));
nor2 add_76_82_g6786 (.a(add_76_82_n_1271), .b(add_76_82_n_1302), .y(n_1645));
nor2 add_76_69_g6787 (.a(add_76_69_n_1024), .b(add_76_69_n_1104), .y(n_1646));
xor2 g6406__6789 (.a(n_1655), .b(n_2618), .y(n_1656));
xor2 add_76_82_g6790 (.a(n_1653), .b(n_1654), .y(n_1655));
xor2 add_76_69_g6791 (.a(n_1651), .b(n_1652), .y(n_1653));
nor2 add_76_82_g6792 (.a(add_76_82_n_1211), .b(add_76_82_n_1299), .y(n_1651));
nor2 add_76_69_g6793 (.a(add_76_69_n_1027), .b(add_76_69_n_1043), .y(n_1652));
nand2 add_76_69_g6794 (.a(add_76_69_n_656), .b(n_2320), .y(n_1654));
nor2 add_76_21_g6795 (.a(n_1661), .b(v0_26_), .y(n_1662));
xor2 g6404__6796 (.a(n_2330), .b(n_1660), .y(n_1661));
nand2 add_76_82_g6799 (.a(add_76_82_n_1291), .b(add_76_82_n_1234), .y(n_1658));
nor2 add_76_82_g6800 (.a(add_76_82_n_839), .b(add_76_82_n_863), .y(n_1660));
nand2 add_76_21_g6801 (.a(n_1661), .b(v0_26_), .y(n_1663));
xor2 add_76_82_g6803 (.a(n_1666), .b(n_1667), .y(n_1668));
xor2 add_76_69_g6804 (.a(n_1664), .b(n_1665), .y(n_1666));
nor2 add_76_82_g6805 (.a(add_76_82_n_1270), .b(add_76_82_n_1285), .y(n_1664));
nor2 add_76_69_g6806 (.a(add_76_69_n_1004), .b(add_76_69_n_1096), .y(n_1665));
nand2 add_76_69_g6807 (.a(add_76_69_n_674), .b(add_76_69_n_655), .y(n_1667));
nand2 g919 (.a(n_1682), .b(n_1690), .y(n_1691));
nand2 g923 (.a(n_1673), .b(n_1681), .y(n_1682));
inv g926 (.a(n_1672), .y(n_1673));
nor2 g927 (.a(n_1670), .b(n_1671), .y(n_1672));
nand2 g933 (.a(add_88_21_n_673), .b(n_2852), .y(n_1670));
nand2 g936 (.a(add_88_21_n_774), .b(n_1782), .y(n_1671));
nor2 g925 (.a(n_1678), .b(n_4371), .y(n_1681));
inv g931 (.a(n_1677), .y(n_1678));
nand2 g932 (.a(n_1674), .b(n_1676), .y(n_1677));
nand2 g937 (.a(n_2126), .b(v1_29_), .y(n_1674));
inv g934 (.a(n_2125), .y(n_1676));
nor2 g920 (.a(n_1687), .b(n_1689), .y(n_1690));
nor2 g921 (.a(n_1670), .b(n_1686), .y(n_1687));
nand2 g922 (.a(add_88_21_n_774), .b(n_1685), .y(n_1686));
nor2 g924 (.a(n_1684), .b(n_1677), .y(n_1685));
nand2 g930 (.a(n_1782), .b(n_1683), .y(n_1684));
inv g928 (.a(n_1688), .y(n_1689));
nand2 g929 (.a(n_4371), .b(v1_r_29_), .y(n_1688));
nand2 g994 (.a(n_1705), .b(n_1709), .y(n_1710));
inv g995 (.a(n_1704), .y(n_1705));
nand2 g996 (.a(n_1702), .b(n_1703), .y(n_1704));
nand2 g997 (.a(n_1700), .b(n_1701), .y(n_1702));
nor2 g998 (.a(add_88_21_n_681), .b(n_1699), .y(n_1700));
inv g1000 (.a(n_1698), .y(n_1699));
nor2 g1001 (.a(add_88_21_n_806), .b(n_4003), .y(n_1698));
nor2 g1009 (.a(add_88_21_n_743), .b(add_88_21_n_773), .y(n_1701));
nand2 g1006 (.a(n_4371), .b(v1_r_31_), .y(n_1703));
nand2 g999 (.a(n_1707), .b(n_4002), .y(n_1709));
nand2 g1005 (.a(n_1706), .b(n_1701), .y(n_1707));
nor2 g1008 (.a(add_88_21_n_681), .b(add_88_21_n_806), .y(n_1706));
nand2 g488 (.a(n_1724), .b(n_1730), .y(n_1731));
mux2 g489 (.a(n_1718), .b(n_1723), .sel(add_88_21_n_731), .y(n_1724));
nand2 g496 (.a(n_1714), .b(n_1683), .y(n_1718));
nand2 g497 (.a(n_1711), .b(n_1713), .y(n_1714));
nand2 g503 (.a(n_1453), .b(v1_25_), .y(n_1711));
inv g504 (.a(n_1712), .y(n_1713));
nor2 g505 (.a(n_1453), .b(v1_25_), .y(n_1712));
nand2 g493 (.a(n_1719), .b(n_1722), .y(n_1723));
nand2 g501 (.a(add_88_21_n_693), .b(add_88_21_n_789), .y(n_1719));
nor2 g494 (.a(n_1721), .b(n_1714), .y(n_1722));
nand2 g498 (.a(add_88_21_n_1119), .b(n_1683), .y(n_1721));
nor2 g490 (.a(n_1725), .b(n_1729), .y(n_1730));
nor2 g491 (.a(n_1719), .b(n_1718), .y(n_1725));
nand2 g492 (.a(n_1727), .b(n_1728), .y(n_1729));
nand2 g495 (.a(n_1726), .b(n_1714), .y(n_1727));
nor2 g500 (.a(add_88_21_n_1119), .b(n_4371), .y(n_1726));
nand2 g499 (.a(n_4371), .b(v1_r_25_), .y(n_1728));
inv g502 (.a(n_1711), .y(n_1732));
inv g560 (.a(n_1755), .y(n_1756));
nor2 g561 (.a(n_1747), .b(n_1754), .y(n_1755));
mux2 g562 (.a(n_1741), .b(n_1746), .sel(add_88_21_n_734), .y(n_1747));
nor2 g563 (.a(n_1733), .b(n_1740), .y(n_1741));
nor2 g577 (.a(n_3284), .b(add_88_21_n_791), .y(n_1733));
nand2 g566 (.a(add_88_21_n_897), .b(n_3442), .y(n_1740));
inv g582 (.a(v1_26_), .y(n_1737));
nor2 g571 (.a(n_1745), .b(n_4371), .y(n_1746));
nor2 g575 (.a(add_88_21_n_1060), .b(n_2118), .y(n_1745));
inv g578 (.a(n_1742), .y(add_88_21_n_1060));
nand2 g579 (.a(n_2119), .b(v1_26_), .y(n_1742));
nand2 g564 (.a(n_1748), .b(n_1753), .y(n_1754));
nand2 g568 (.a(n_1733), .b(n_1746), .y(n_1748));
nor2 g565 (.a(n_1750), .b(n_1752), .y(n_1753));
nor2 g567 (.a(add_88_21_n_897), .b(n_1749), .y(n_1750));
inv g570 (.a(n_1746), .y(n_1749));
inv g572 (.a(n_1751), .y(n_1752));
nand2 g573 (.a(n_4371), .b(v1_r_26_), .y(n_1751));
inv g767 (.a(n_1757), .y(n_1758));
nor2 g768 (.a(add_88_21_n_803), .b(n_3284), .y(n_1757));
nor2 g757 (.a(n_1766), .b(n_4371), .y(n_1769));
inv g763 (.a(n_1765), .y(n_1766));
nand2 g764 (.a(n_1762), .b(n_1764), .y(n_1765));
nand2 g769 (.a(n_2202), .b(v1_27_), .y(n_1762));
inv g765 (.a(n_2201), .y(n_1764));
nor2 g752 (.a(n_1773), .b(n_1775), .y(n_1776));
nor2 g753 (.a(n_2499), .b(n_1772), .y(n_1773));
nand2 g755 (.a(add_88_21_n_787), .b(n_1771), .y(n_1772));
nor2 g758 (.a(n_1765), .b(n_4371), .y(n_1771));
inv g761 (.a(n_1774), .y(n_1775));
nand2 g762 (.a(n_4371), .b(v1_r_27_), .y(n_1774));
nand2 g6811 (.a(add_88_21_n_810), .b(add_88_21_n_693), .y(n_1779));
nand2 g6812 (.a(n_1785), .b(n_1683), .y(n_1789));
nand2 g6813 (.a(n_1782), .b(n_2854), .y(n_1785));
nand2 g6814 (.a(n_2131), .b(v1_28_), .y(n_1782));
inv g6817 (.a(n_4371), .y(n_1683));
nand2 g747 (.a(n_1795), .b(n_1796), .y(n_1797));
nand2 g748 (.a(n_1791), .b(n_1794), .y(n_1795));
inv g6820 (.a(n_2507), .y(n_1791));
nor2 g750 (.a(add_88_21_n_797), .b(n_1793), .y(n_1794));
nand2 g6821 (.a(n_1792), .b(n_1683), .y(n_1793));
inv g6822 (.a(n_1785), .y(n_1792));
nand2 g6823 (.a(n_4371), .b(v1_r_28_), .y(n_1796));
nor2 g6828 (.a(n_1803), .b(n_1807), .y(n_1808));
nand2 g6829 (.a(add_88_21_n_868), .b(n_1683), .y(n_1803));
inv g944 (.a(ps_0_), .y(n_1800));
nand2 g6830 (.a(n_1804), .b(n_1806), .y(n_1807));
nand2 g941 (.a(n_2998), .b(v1_30_), .y(n_1804));
inv g6831 (.a(n_1805), .y(n_1806));
nor2 g939 (.a(n_2998), .b(v1_30_), .y(n_1805));
nand2 g6832 (.a(add_88_21_n_741), .b(add_88_21_n_764), .y(n_1810));
inv g6833 (.a(n_1812), .y(n_1813));
nand2 g6834 (.a(n_4371), .b(v1_r_30_), .y(n_1812));
nand2 g6835 (.a(n_1817), .b(n_1819), .y(n_1820));
inv g6836 (.a(n_1816), .y(n_1817));
nor2 g6837 (.a(n_1810), .b(n_1815), .y(n_1816));
nand2 g940 (.a(add_88_21_n_688), .b(add_88_21_n_868), .y(n_1815));
nor2 g6838 (.a(n_1818), .b(n_4371), .y(n_1819));
inv g6839 (.a(n_1807), .y(n_1818));
nor2 g597 (.a(add_76_21_n_1238), .b(n_1322), .y(n_1827));
nor2 g293 (.a(n_2683), .b(n_1845), .y(n_1846));
nand2 g297 (.a(n_2905), .b(n_1844), .y(n_1845));
inv g301 (.a(n_1843), .y(n_1844));
nor2 g302 (.a(n_1842), .b(sum_4_), .y(n_1843));
inv g309 (.a(n_1841), .y(n_1842));
nor2 g310 (.a(n_502), .b(n_501), .y(n_1841));
inv g294 (.a(n_1849), .y(n_1850));
nor2 g295 (.a(n_2914), .b(n_1848), .y(n_1849));
nand2 g312 (.a(n_1861), .b(n_2901), .y(n_1848));
nand2 g623 (.a(n_1862), .b(n_1867), .y(n_1868));
nand2 g625 (.a(n_3125), .b(n_1861), .y(n_1862));
nand2 g630 (.a(n_1860), .b(sum_1_), .y(n_1861));
inv g632 (.a(n_1859), .y(n_1860));
nor2 g633 (.a(n_493), .b(n_492), .y(n_1859));
nor2 g628 (.a(n_2681), .b(n_1866), .y(n_1867));
nor2 g629 (.a(n_1860), .b(sum_1_), .y(n_1866));
inv g626 (.a(n_1869), .y(n_1870));
nor2 g627 (.a(n_3125), .b(n_1866), .y(n_1869));
nor2 g6844 (.a(n_4290), .b(n_1881), .y(n_1882));
nand2 g6850 (.a(n_4499), .b(add_76_21_n_1209), .y(n_1881));
inv g600 (.a(n_3881), .y(add_76_21_n_1209));
nor2 g6852 (.a(n_1887), .b(n_1889), .y(n_1890));
nor2 g583 (.a(n_1884), .b(n_1886), .y(n_1887));
inv g602 (.a(n_3664), .y(n_1884));
nand2 g6853 (.a(n_1885), .b(n_1881), .y(n_1886));
nor2 g6854 (.a(n_1985), .b(n_4291), .y(n_1885));
nor2 g6855 (.a(n_4289), .b(n_1888), .y(n_1889));
inv g6856 (.a(n_1881), .y(n_1888));
inv g6858 (.a(n_1886), .y(n_1892));
nand2 g6859 (.a(n_4289), .b(n_1894), .y(n_1895));
nor2 g6860 (.a(n_1885), .b(n_1881), .y(n_1894));
inv g398 (.a(n_1905), .y(n_1906));
nor2 g399 (.a(add_88_69_n_1648), .b(n_1904), .y(n_1905));
nor2 g401 (.a(n_2586), .b(n_2033), .y(n_1904));
nand2 g409 (.a(n_3525), .b(n_1224), .y(n_1910));
nand2 g402 (.a(n_1916), .b(n_1918), .y(n_1919));
nor2 g403 (.a(n_1914), .b(n_1915), .y(n_1916));
nor2 g410 (.a(add_88_69_n_1717), .b(add_88_69_n_1648), .y(n_1914));
inv g408 (.a(n_1910), .y(n_1915));
nand2 g404 (.a(n_2039), .b(n_1917), .y(n_1918));
nor2 g407 (.a(add_88_69_n_1668), .b(add_88_69_n_1648), .y(n_1917));
nor2 g1074 (.a(n_1922), .b(n_2310), .y(n_1924));
inv g1080 (.a(n_1921), .y(n_1922));
nand2 g1081 (.a(n_2311), .b(v0_25_), .y(n_1921));
nor2 g1069 (.a(n_1928), .b(n_1929), .y(n_1930));
nand2 g1073 (.a(n_1924), .b(n_1927), .y(n_1928));
nand2 g1077 (.a(n_1656), .b(v0_24_), .y(n_1927));
inv g1084 (.a(n_1605), .y(n_1929));
nor2 g1071 (.a(n_1924), .b(n_1927), .y(n_1931));
nand2 g1067 (.a(n_3710), .b(n_1935), .y(n_1936));
inv g1072 (.a(n_1928), .y(n_1935));
nor2 g1061 (.a(n_3955), .b(n_3710), .y(n_1941));
inv g1076 (.a(n_1927), .y(n_1946));
nor2 g740 (.a(n_1950), .b(n_1955), .y(n_1956));
nand2 g6861 (.a(n_3941), .b(add_76_21_n_932), .y(n_1950));
inv g6862 (.a(n_1948), .y(add_76_21_n_932));
nand2 g6863 (.a(add_76_21_n_981), .b(add_76_21_n_1018), .y(n_1948));
nand2 g743 (.a(add_76_21_n_950), .b(n_1954), .y(n_1955));
nor2 g6864 (.a(n_1952), .b(n_3010), .y(n_1954));
inv g6865 (.a(n_3011), .y(n_1952));
nor2 g741 (.a(n_3954), .b(n_1963), .y(n_1964));
nor2 g6869 (.a(n_3710), .b(add_76_21_n_950), .y(n_1959));
nand2 g6871 (.a(add_76_21_n_1016), .b(n_1962), .y(n_1963));
inv g6873 (.a(n_1954), .y(n_1962));
nor2 g737 (.a(n_1968), .b(n_1970), .y(n_1971));
nor2 g742 (.a(n_1966), .b(n_1967), .y(n_1968));
nand2 g6874 (.a(n_3941), .b(n_3710), .y(n_1966));
nand2 g6875 (.a(add_76_21_n_932), .b(n_1954), .y(n_1967));
mux2 g739 (.a(n_1962), .b(n_1969), .sel(n_1948), .y(n_1970));
nor2 g6876 (.a(add_76_21_n_1016), .b(n_1962), .y(n_1969));
nor2 g334 (.a(n_3660), .b(n_3709), .y(n_1983));
nand2 g341 (.a(n_1977), .b(n_4292), .y(n_1980));
nor2 g346 (.a(n_4502), .b(n_4291), .y(n_1977));
mux2 g339 (.a(n_1984), .b(n_1985), .sel(n_1986), .y(n_1987));
inv g343 (.a(n_4292), .y(n_1984));
nor2 g342 (.a(n_3869), .b(v0_16_), .y(n_1985));
inv g345 (.a(n_1977), .y(n_1986));
nand2 g338 (.a(n_3709), .b(n_1989), .y(n_1990));
nor2 g340 (.a(n_1977), .b(n_1985), .y(n_1989));
nand2 g335 (.a(n_3664), .b(n_1989), .y(n_1991));
xor2 g785 (.a(n_1996), .b(n_1997), .y(n_1998));
nor2 g791 (.a(add_76_21_n_893), .b(add_76_21_n_861), .y(n_1996));
nand2 g788 (.a(n_1400), .b(add_76_21_n_1181), .y(n_1997));
xor2 g779 (.a(n_2005), .b(n_2085), .y(n_2007));
xor2 g784 (.a(n_2003), .b(n_2004), .y(n_2005));
nor2 g792 (.a(add_76_21_n_940), .b(add_76_21_n_863), .y(n_2003));
nand2 g790 (.a(n_1421), .b(add_76_21_n_1254), .y(n_2004));
nor2 g645 (.a(n_2014), .b(n_3694), .y(n_2017));
inv g648 (.a(n_3692), .y(n_2014));
nand2 g642 (.a(n_2018), .b(n_2019), .y(n_2020));
nand2 g652 (.a(n_3701), .b(v0_8_), .y(n_2018));
nand2 g647 (.a(n_3693), .b(v0_9_), .y(n_2019));
nor2 g221 (.a(n_2028), .b(n_2037), .y(n_2038));
nor2 g226 (.a(n_2025), .b(n_2027), .y(n_2028));
nor2 g232 (.a(n_3967), .b(add_88_69_n_1699), .y(n_2025));
inv g233 (.a(n_2026), .y(n_2027));
nor2 g234 (.a(add_88_69_n_1668), .b(n_1906), .y(n_2026));
nand2 g222 (.a(n_2030), .b(n_2036), .y(n_2037));
inv g229 (.a(n_2029), .y(n_2030));
nor2 g230 (.a(add_88_69_n_1717), .b(n_1906), .y(n_2029));
nor2 g223 (.a(n_2031), .b(n_2035), .y(n_2036));
nor2 g235 (.a(n_1910), .b(n_1904), .y(n_2031));
inv g224 (.a(n_2034), .y(n_2035));
nand2 g225 (.a(n_2586), .b(n_2033), .y(n_2034));
xor2 g227 (.a(add_76_21_n_800), .b(add_76_21_n_1122), .y(n_2033));
inv g231 (.a(n_2025), .y(n_2039));
mux2 g381 (.a(n_2042), .b(n_2043), .sel(n_4058), .y(n_2049));
nor2 g387 (.a(n_2041), .b(v0_29_), .y(n_2042));
inv g390 (.a(n_3984), .y(n_2041));
nor2 g386 (.a(n_3984), .b(v0_29_), .y(n_2043));
nor2 g389 (.a(add_76_69_n_665), .b(add_76_69_n_651), .y(n_2044));
nand2 g388 (.a(add_76_69_n_1012), .b(add_76_69_n_1082), .y(n_2045));
nor2 g6878 (.a(n_2054), .b(n_2057), .y(n_2058));
nand2 g6879 (.a(n_3744), .b(n_3761), .y(n_2054));
nand2 g6880 (.a(n_3779), .b(n_3796), .y(n_2057));
inv g6883 (.a(n_2058), .y(n_2060));
nand2 g6885 (.a(n_2068), .b(n_2074), .y(n_2075));
nand2 g6886 (.a(n_2063), .b(n_2067), .y(n_2068));
inv g6887 (.a(n_2062), .y(n_2063));
nor2 g593 (.a(n_2058), .b(sum_0_), .y(n_2062));
nand2 g6888 (.a(n_2065), .b(n_2066), .y(n_2067));
inv g6889 (.a(n_2064), .y(n_2065));
nor2 g6890 (.a(n_3821), .b(n_3830), .y(n_2064));
xor2 g6891 (.a(sum_0_), .b(sum_1_), .y(n_2066));
nor2 g6892 (.a(n_2069), .b(n_2073), .y(n_2074));
nor2 g6893 (.a(n_2065), .b(n_2066), .y(n_2069));
nor2 g6894 (.a(n_2072), .b(n_457), .y(n_2073));
inv g6895 (.a(n_2071), .y(n_2072));
nor2 g6896 (.a(n_3839), .b(n_2070), .y(n_2071));
xor2 g591 (.a(inc_add_77_23_n_527), .b(inc_add_77_23_n_566), .y(n_2070));
nand2 g6897 (.a(n_2077), .b(n_2067), .y(n_2078));
nand2 g6898 (.a(n_2062), .b(n_2076), .y(n_2077));
inv g6899 (.a(n_2069), .y(n_2076));
inv g594 (.a(n_2079), .y(n_2080));
nor2 g6900 (.a(n_3839), .b(n_457), .y(n_2079));
nand2 g853 (.a(n_1550), .b(add_76_21_n_1277), .y(n_2085));
mux2 g841 (.a(n_2091), .b(n_2092), .sel(n_4059), .y(n_2096));
nor2 g844 (.a(n_2089), .b(n_4306), .y(n_2091));
inv g854 (.a(n_3493), .y(n_2089));
nor2 g843 (.a(n_3493), .b(n_4306), .y(n_2092));
nand2 g1216 (.a(n_2105), .b(n_2109), .y(n_2110));
nand2 g1219 (.a(n_2101), .b(n_2104), .y(n_2105));
nor2 g1221 (.a(n_2099), .b(n_2100), .y(n_2101));
nor2 g1227 (.a(n_3599), .b(add_88_69_n_1491), .y(n_2099));
nand2 g1226 (.a(add_88_69_n_1437), .b(add_88_69_n_1717), .y(n_2100));
nand2 g1220 (.a(n_2102), .b(n_2103), .y(n_2104));
nor2 g1223 (.a(add_88_69_n_1408), .b(add_88_69_n_1491), .y(n_2102));
nand2 g1225 (.a(add_88_69_n_1292), .b(add_88_69_n_1322), .y(n_2103));
inv g1217 (.a(n_2108), .y(n_2109));
xor2 g1218 (.a(n_2106), .b(n_2107), .y(n_2108));
xor2 g1222 (.a(add_88_82_n_1917), .b(add_88_82_n_2143), .y(n_2106));
nor2 g1224 (.a(n_1915), .b(add_88_69_n_1648), .y(n_2107));
nand2 g1213 (.a(n_2112), .b(n_2101), .y(n_2113));
inv g1214 (.a(n_2111), .y(n_2112));
nand2 g1215 (.a(n_2104), .b(n_2108), .y(n_2111));
mux2 g57 (.a(n_2116), .b(n_2117), .sel(n_1348), .y(n_2118));
nor2 g60 (.a(n_2115), .b(v1_26_), .y(n_2116));
inv g61 (.a(n_1347), .y(n_2115));
nor2 g59 (.a(n_1347), .b(v1_26_), .y(n_2117));
xor2 g58 (.a(n_1348), .b(n_1347), .y(n_2119));
xor2 g41 (.a(add_88_69_n_1243), .b(n_2120), .y(n_2121));
xor2 g42 (.a(n_825), .b(n_3966), .y(n_2120));
mux2 g72 (.a(n_2123), .b(n_2124), .sel(n_1362), .y(n_2125));
nor2 g75 (.a(n_2122), .b(v1_29_), .y(n_2123));
inv g76 (.a(n_1361), .y(n_2122));
nor2 g74 (.a(n_1361), .b(v1_29_), .y(n_2124));
xor2 g73 (.a(n_1362), .b(n_1361), .y(n_2126));
xor2 g6905 (.a(n_4019), .b(n_4022), .y(n_2131));
nand2 g25 (.a(n_2133), .b(n_2134), .y(n_2135));
nor2 g27 (.a(n_3891), .b(n_1316), .y(n_2133));
inv g28 (.a(n_2846), .y(n_1316));
inv g29 (.a(add_88_21_n_895), .y(n_2134));
nor2 g26 (.a(add_88_21_n_895), .b(n_3891), .y(n_2136));
inv g89 (.a(n_2137), .y(n_2138));
nor2 g90 (.a(add_88_21_n_1006), .b(n_4371), .y(n_2137));
nand2 g92 (.a(add_88_21_n_1006), .b(n_1683), .y(n_2140));
nand2 g91 (.a(n_4371), .b(v1_r_17_), .y(n_2142));
inv g6908 (.a(n_2144), .y(n_2145));
nor2 g6909 (.a(add_88_21_n_1002), .b(n_4371), .y(n_2144));
nand2 g6910 (.a(add_88_21_n_1002), .b(n_1683), .y(n_2147));
nand2 g6912 (.a(n_4371), .b(v1_r_18_), .y(n_2149));
inv g6915 (.a(n_2151), .y(n_2152));
nor2 g6916 (.a(add_88_21_n_996), .b(n_4371), .y(n_2151));
nand2 g6917 (.a(add_88_21_n_996), .b(n_1683), .y(n_2154));
nand2 g6919 (.a(n_4371), .b(v1_r_19_), .y(n_2156));
inv g6922 (.a(n_2158), .y(n_2159));
nor2 g6923 (.a(add_88_21_n_1003), .b(n_4371), .y(n_2158));
nand2 g6924 (.a(add_88_21_n_1003), .b(n_1683), .y(n_2161));
nand2 g6926 (.a(n_4371), .b(v1_r_20_), .y(n_2163));
inv g6929 (.a(n_2165), .y(n_2166));
nor2 g6930 (.a(add_88_21_n_989), .b(n_4371), .y(n_2165));
nand2 g6931 (.a(add_88_21_n_989), .b(n_1683), .y(n_2168));
nand2 g6933 (.a(n_4371), .b(v1_r_21_), .y(n_2170));
inv g6936 (.a(n_2172), .y(n_2173));
nor2 g6937 (.a(add_88_21_n_980), .b(n_4371), .y(n_2172));
nand2 g6938 (.a(add_88_21_n_980), .b(n_1683), .y(n_2175));
nand2 g6940 (.a(n_4371), .b(v1_r_22_), .y(n_2177));
nor2 g6944 (.a(add_88_21_n_991), .b(n_4371), .y(n_2179));
nand2 g6945 (.a(add_88_21_n_991), .b(n_1683), .y(n_2182));
nand2 g6947 (.a(n_4371), .b(v1_r_23_), .y(n_2184));
inv g6950 (.a(n_2186), .y(n_2187));
nor2 g6951 (.a(add_88_21_n_1020), .b(n_4371), .y(n_2186));
nand2 g6952 (.a(add_88_21_n_1020), .b(n_1683), .y(n_2189));
nand2 g6954 (.a(n_4371), .b(v1_r_24_), .y(n_2191));
xor2 g6955 (.a(n_2193), .b(add_76_21_n_804), .y(n_2194));
xor2 g6956 (.a(n_2961), .b(add_76_21_n_1121), .y(n_2193));
xor2 g6957 (.a(add_76_21_n_804), .b(add_76_21_n_1121), .y(n_2195));
xor2 g31 (.a(n_2103), .b(n_2196), .y(n_2197));
xor2 g32 (.a(add_88_69_n_1612), .b(n_801), .y(n_2196));
nor2 g24 (.a(n_2199), .b(n_2200), .y(n_2201));
nand2 g6958 (.a(n_2113), .b(n_2198), .y(n_2199));
inv g6959 (.a(v1_27_), .y(n_2198));
inv g6960 (.a(n_2110), .y(n_2200));
nand2 g6961 (.a(n_2110), .b(n_2113), .y(n_2202));
inv g280 (.a(n_3956), .y(n_2211));
nor2 g284 (.a(n_2520), .b(n_2096), .y(n_2204));
nand2 g95 (.a(n_2215), .b(n_2218), .y(n_2219));
nor2 g98 (.a(n_2213), .b(n_2214), .y(n_2215));
nor2 g102 (.a(add_76_82_n_896), .b(n_2212), .y(n_2213));
inv g103 (.a(add_76_82_n_981), .y(n_2212));
inv g104 (.a(add_76_82_n_901), .y(n_2214));
nand2 g97 (.a(n_2362), .b(n_2217), .y(n_2218));
inv g99 (.a(n_2216), .y(n_2217));
nand2 g100 (.a(add_76_82_n_981), .b(n_2579), .y(n_2216));
nand2 g6962 (.a(n_2227), .b(n_2229), .y(n_2230));
nand2 g507 (.a(n_2225), .b(n_2226), .y(n_2227));
nand2 g508 (.a(n_2223), .b(n_2224), .y(n_2225));
inv g510 (.a(n_2222), .y(n_2223));
nor2 g511 (.a(add_76_69_n_664), .b(add_76_69_n_800), .y(n_2222));
inv g512 (.a(add_76_69_n_707), .y(n_2224));
xor2 g6963 (.a(n_1633), .b(add_76_69_n_948), .y(n_2226));
nand2 g6964 (.a(n_2223), .b(n_2228), .y(n_2229));
nor2 g6965 (.a(add_76_69_n_707), .b(n_2226), .y(n_2228));
nor2 g6968 (.a(add_76_82_n_896), .b(n_2231), .y(n_2232));
inv g6969 (.a(add_76_82_n_1075), .y(n_2231));
inv g6970 (.a(add_76_82_n_951), .y(n_2233));
nand2 g6971 (.a(n_2362), .b(n_2236), .y(n_2237));
inv g6972 (.a(n_2235), .y(n_2236));
nand2 g6973 (.a(n_2579), .b(add_76_82_n_1075), .y(n_2235));
nor2 g454 (.a(n_2247), .b(n_2250), .y(n_2251));
nor2 g457 (.a(n_3843), .b(n_2246), .y(n_2247));
nand2 g461 (.a(n_1528), .b(add_76_69_n_1036), .y(n_2246));
mux2 g456 (.a(add_76_69_n_1090), .b(add_76_69_n_1035), .sel(n_1528), .y(n_2250));
inv g464 (.a(add_76_69_n_1036), .y(add_76_69_n_1035));
nor2 g455 (.a(n_2254), .b(n_2255), .y(n_2256));
nor2 g459 (.a(n_2566), .b(n_4558), .y(n_2254));
nor2 g458 (.a(n_2565), .b(n_4558), .y(n_2255));
nand2 g143 (.a(n_2261), .b(add_76_82_n_1293), .y(n_2262));
nand2 g147 (.a(n_2581), .b(add_76_82_n_954), .y(n_2261));
nand2 g429 (.a(n_2272), .b(n_2276), .y(n_2277));
nand2 g433 (.a(n_2601), .b(n_2271), .y(n_2272));
inv g435 (.a(n_2270), .y(n_2271));
nor2 g436 (.a(n_2269), .b(add_76_82_n_911), .y(n_2270));
nor2 g437 (.a(n_3648), .b(add_76_82_n_1022), .y(n_2269));
inv g431 (.a(n_2275), .y(n_2276));
nor2 g432 (.a(n_2274), .b(n_2269), .y(n_2275));
nand2 g434 (.a(n_2602), .b(n_2273), .y(n_2274));
nor2 g438 (.a(add_76_82_n_911), .b(v0_15_), .y(n_2273));
xor2 g430 (.a(n_2270), .b(n_2602), .y(n_2278));
nand2 g6976 (.a(n_2283), .b(n_2287), .y(n_2288));
nand2 g6977 (.a(n_2279), .b(n_2282), .y(n_2283));
nor2 g6978 (.a(n_1473), .b(v0_14_), .y(n_2279));
inv g6979 (.a(n_2281), .y(n_2282));
nor2 g6980 (.a(n_2280), .b(add_76_82_n_903), .y(n_2281));
nor2 g6981 (.a(n_3648), .b(add_76_82_n_996), .y(n_2280));
inv g6982 (.a(n_2286), .y(n_2287));
nor2 g6983 (.a(n_2285), .b(n_2280), .y(n_2286));
nand2 g6984 (.a(n_1473), .b(n_2284), .y(n_2285));
nor2 g6985 (.a(add_76_82_n_903), .b(v0_14_), .y(n_2284));
xor2 g6986 (.a(n_2281), .b(n_1473), .y(n_2289));
nand2 g6987 (.a(n_2294), .b(n_2298), .y(n_2299));
nand2 g6988 (.a(n_2291), .b(n_2293), .y(n_2294));
nor2 g414 (.a(n_2290), .b(v0_13_), .y(n_2291));
inv g417 (.a(n_1447), .y(n_2290));
nand2 g411 (.a(n_2292), .b(add_76_82_n_902), .y(n_2293));
nand2 g413 (.a(n_2362), .b(add_76_82_n_986), .y(n_2292));
nand2 g6989 (.a(n_2297), .b(n_2292), .y(n_2298));
nor2 g412 (.a(n_1447), .b(n_2296), .y(n_2297));
nand2 g415 (.a(add_76_82_n_902), .b(n_2295), .y(n_2296));
inv g416 (.a(v0_13_), .y(n_2295));
xor2 g6990 (.a(n_2293), .b(n_1447), .y(n_2300));
nand2 g6991 (.a(n_2305), .b(n_2309), .y(n_2310));
nand2 g6992 (.a(n_2630), .b(n_2304), .y(n_2305));
nand2 g6995 (.a(n_2303), .b(n_2658), .y(n_2304));
nand2 g6996 (.a(n_3866), .b(add_76_82_n_946), .y(n_2303));
nand2 g6997 (.a(n_2308), .b(n_2303), .y(n_2309));
nor2 g6998 (.a(n_2649), .b(n_2657), .y(n_2308));
xor2 g7001 (.a(n_2304), .b(n_2649), .y(n_2311));
inv g119 (.a(n_2317), .y(n_2318));
nor2 g120 (.a(n_2313), .b(n_2316), .y(n_2317));
nand2 g121 (.a(n_2312), .b(add_76_69_n_837), .y(n_2313));
nand2 g125 (.a(add_76_69_n_767), .b(add_76_69_n_901), .y(n_2312));
nor2 g124 (.a(add_76_69_n_744), .b(n_2315), .y(n_2316));
nand2 g127 (.a(n_2314), .b(add_76_69_n_901), .y(n_2315));
inv g128 (.a(add_76_69_n_833), .y(n_2314));
inv g122 (.a(n_2320), .y(n_2321));
nor2 g123 (.a(n_2319), .b(add_76_69_n_767), .y(n_2320));
nor2 g126 (.a(add_76_69_n_744), .b(add_76_69_n_833), .y(n_2319));
nand2 g7002 (.a(n_2327), .b(n_2329), .y(n_2330));
nand2 g7003 (.a(n_2325), .b(n_2326), .y(n_2327));
nand2 g7004 (.a(n_2323), .b(n_2317), .y(n_2325));
inv g7005 (.a(n_2322), .y(n_2323));
nor2 g7006 (.a(add_76_69_n_664), .b(add_76_69_n_757), .y(n_2322));
xor2 g7008 (.a(n_1658), .b(add_76_69_n_935), .y(n_2326));
nand2 g7009 (.a(n_2328), .b(n_2323), .y(n_2329));
nor2 g7010 (.a(n_2318), .b(n_2326), .y(n_2328));
nand2 g7011 (.a(n_2335), .b(n_2339), .y(n_2340));
nand2 g7012 (.a(n_2331), .b(n_2334), .y(n_2335));
nor2 g421 (.a(n_1479), .b(v0_12_), .y(n_2331));
inv g7013 (.a(n_2333), .y(n_2334));
nor2 g418 (.a(n_2332), .b(add_76_82_n_938), .y(n_2333));
nor2 g419 (.a(n_3648), .b(n_2578), .y(n_2332));
inv g7014 (.a(n_2338), .y(n_2339));
nor2 g7015 (.a(n_2337), .b(n_2332), .y(n_2338));
nand2 g7016 (.a(n_1479), .b(n_2336), .y(n_2337));
nor2 g420 (.a(add_76_82_n_938), .b(v0_12_), .y(n_2336));
xor2 g7017 (.a(n_2333), .b(n_1479), .y(n_2341));
nand2 g7019 (.a(n_2741), .b(n_3645), .y(n_2346));
nor2 g7027 (.a(add_76_82_n_948), .b(v0_11_), .y(n_2347));
xor2 g7028 (.a(n_3646), .b(n_3652), .y(n_2352));
nand2 g7029 (.a(add_76_82_n_954), .b(add_76_82_n_1091), .y(n_2353));
nand2 g7030 (.a(n_2807), .b(add_76_82_n_1091), .y(n_2356));
inv g116 (.a(n_3648), .y(n_2362));
nand2 g109 (.a(n_2366), .b(n_3909), .y(n_2370));
nor2 g111 (.a(n_2364), .b(n_2365), .y(n_2366));
nor2 g7033 (.a(n_2363), .b(add_76_82_n_1208), .y(n_2364));
inv g7034 (.a(add_76_82_n_954), .y(n_2363));
inv g7035 (.a(add_76_82_n_1276), .y(n_2365));
xor2 g7039 (.a(n_874), .b(add_76_82_n_1148), .y(n_2373));
nand2 g291 (.a(n_2387), .b(n_2390), .y(n_2391));
nor2 g7041 (.a(n_2379), .b(n_3452), .y(n_2387));
nor2 g7042 (.a(n_3284), .b(n_2378), .y(n_2379));
inv g7043 (.a(n_2377), .y(n_2378));
nor2 g7044 (.a(n_2138), .b(add_88_21_n_1123), .y(n_2377));
nor2 g7047 (.a(n_2138), .b(add_88_21_n_1126), .y(n_2380));
nor2 g7050 (.a(n_2140), .b(add_88_21_n_1122), .y(n_2384));
nand2 g7052 (.a(n_3284), .b(n_2389), .y(n_2390));
nor2 g7053 (.a(n_2140), .b(n_2388), .y(n_2389));
inv g7054 (.a(add_88_21_n_1126), .y(n_2388));
nand2 g7055 (.a(n_2402), .b(n_2405), .y(n_2406));
nor2 g7056 (.a(n_2394), .b(n_2401), .y(n_2402));
nor2 g7057 (.a(add_88_21_n_693), .b(n_2393), .y(n_2394));
nand2 g7058 (.a(n_2392), .b(add_88_21_n_872), .y(n_2393));
inv g315 (.a(n_2147), .y(n_2392));
nand2 g7059 (.a(n_2397), .b(n_2400), .y(n_2401));
nor2 g7060 (.a(n_2395), .b(n_2396), .y(n_2397));
nor2 g7061 (.a(n_2145), .b(add_88_21_n_872), .y(n_2395));
inv g316 (.a(n_2149), .y(n_2396));
nand2 g308 (.a(n_2392), .b(n_2399), .y(n_2400));
nor2 g7062 (.a(add_88_21_n_873), .b(add_88_21_n_924), .y(n_2399));
nand2 g7063 (.a(add_88_21_n_693), .b(n_2404), .y(n_2405));
nor2 g7064 (.a(n_2145), .b(n_2403), .y(n_2404));
inv g314 (.a(add_88_21_n_924), .y(n_2403));
nand2 g7065 (.a(n_2418), .b(n_2420), .y(n_2421));
nor2 g7066 (.a(n_2409), .b(n_2417), .y(n_2418));
nor2 g7067 (.a(n_3284), .b(n_2408), .y(n_2409));
inv g320 (.a(n_2407), .y(n_2408));
nor2 g321 (.a(n_2154), .b(add_88_21_n_906), .y(n_2407));
inv g7068 (.a(n_2416), .y(n_2417));
nor2 g7069 (.a(n_2412), .b(n_2415), .y(n_2416));
nand2 g318 (.a(n_2411), .b(n_2156), .y(n_2412));
nand2 g323 (.a(add_88_21_n_793), .b(n_2410), .y(n_2411));
inv g324 (.a(n_2154), .y(n_2410));
nor2 g7070 (.a(n_2414), .b(add_88_21_n_793), .y(n_2415));
nand2 g322 (.a(n_2151), .b(add_88_21_n_906), .y(n_2414));
nand2 g7071 (.a(n_3284), .b(n_2419), .y(n_2420));
nor2 g319 (.a(add_88_21_n_793), .b(n_2152), .y(n_2419));
nand2 g7072 (.a(n_2425), .b(n_2432), .y(n_2433));
inv g7073 (.a(n_2424), .y(n_2425));
mux2 g7074 (.a(n_2422), .b(n_2423), .sel(n_3284), .y(n_2424));
nor2 g7075 (.a(add_88_21_n_778), .b(n_2159), .y(n_2422));
nor2 g7076 (.a(n_2161), .b(add_88_21_n_882), .y(n_2423));
nor2 g7077 (.a(n_2428), .b(n_2431), .y(n_2432));
nand2 g7078 (.a(n_2427), .b(n_2163), .y(n_2428));
nand2 g7079 (.a(add_88_21_n_778), .b(n_2426), .y(n_2427));
inv g7080 (.a(n_2161), .y(n_2426));
nor2 g7081 (.a(add_88_21_n_778), .b(n_2430), .y(n_2431));
nand2 g7082 (.a(add_88_21_n_882), .b(n_2158), .y(n_2430));
nand2 g373 (.a(n_2440), .b(n_2447), .y(n_2448));
nor2 g376 (.a(n_2436), .b(n_2439), .y(n_2440));
nor2 g378 (.a(n_2435), .b(add_88_21_n_693), .y(n_2436));
nand2 g7084 (.a(add_88_21_n_749), .b(n_2434), .y(n_2435));
inv g7085 (.a(n_2168), .y(n_2434));
nand2 g380 (.a(n_2438), .b(n_2170), .y(n_2439));
inv g7086 (.a(n_2437), .y(n_2438));
nor2 g7087 (.a(add_88_21_n_749), .b(n_2166), .y(n_2437));
inv g374 (.a(n_2446), .y(n_2447));
nand2 g375 (.a(n_2443), .b(n_2445), .y(n_2446));
nand2 g379 (.a(add_88_21_n_693), .b(n_2442), .y(n_2443));
nor2 g7088 (.a(n_2441), .b(n_2166), .y(n_2442));
inv g7089 (.a(add_88_21_n_820), .y(n_2441));
nand2 g377 (.a(add_88_21_n_749), .b(n_2444), .y(n_2445));
nor2 g7090 (.a(add_88_21_n_820), .b(n_2168), .y(n_2444));
nand2 g7091 (.a(n_2457), .b(n_2462), .y(n_2463));
nor2 g7092 (.a(n_2451), .b(n_2456), .y(n_2457));
inv g7093 (.a(n_2450), .y(n_2451));
nand2 g7094 (.a(n_2449), .b(n_3284), .y(n_2450));
nor2 g7095 (.a(add_88_21_n_750), .b(n_2173), .y(n_2449));
nand2 g7096 (.a(n_2455), .b(n_2177), .y(n_2456));
nand2 g7097 (.a(n_2452), .b(n_2454), .y(n_2455));
inv g7098 (.a(add_88_21_n_750), .y(n_2452));
nor2 g7099 (.a(n_2453), .b(n_2173), .y(n_2454));
inv g7100 (.a(add_88_21_n_828), .y(n_2453));
nor2 g7101 (.a(n_2460), .b(n_2461), .y(n_2462));
nor2 g7102 (.a(n_3284), .b(n_2459), .y(n_2460));
inv g7103 (.a(n_2458), .y(n_2459));
nor2 g7104 (.a(add_88_21_n_828), .b(n_2175), .y(n_2458));
nor2 g7105 (.a(n_2452), .b(n_2175), .y(n_2461));
nand2 g7106 (.a(n_2472), .b(n_2477), .y(n_2478));
nor2 g7107 (.a(n_3233), .b(n_2471), .y(n_2472));
nand2 g7111 (.a(n_2470), .b(n_2184), .y(n_2471));
nand2 g7112 (.a(n_2467), .b(n_3436), .y(n_2470));
inv g7113 (.a(add_88_21_n_758), .y(n_2467));
nor2 g7116 (.a(n_2475), .b(n_2476), .y(n_2477));
nor2 g7117 (.a(n_3284), .b(n_2474), .y(n_2475));
inv g7118 (.a(n_2473), .y(n_2474));
nor2 g7119 (.a(add_88_21_n_860), .b(n_2182), .y(n_2473));
nor2 g7120 (.a(n_2467), .b(n_2182), .y(n_2476));
nand2 g7121 (.a(n_2485), .b(n_2492), .y(n_2493));
nor2 g7122 (.a(n_2481), .b(n_2484), .y(n_2485));
nor2 g7123 (.a(n_2480), .b(add_88_21_n_693), .y(n_2481));
nand2 g7124 (.a(add_88_21_n_746), .b(n_2479), .y(n_2480));
inv g7125 (.a(n_2189), .y(n_2479));
nand2 g7126 (.a(n_2483), .b(n_2191), .y(n_2484));
inv g7127 (.a(n_2482), .y(n_2483));
nor2 g7128 (.a(add_88_21_n_746), .b(n_2187), .y(n_2482));
inv g7129 (.a(n_2491), .y(n_2492));
nand2 g7130 (.a(n_2488), .b(n_2490), .y(n_2491));
nand2 g7131 (.a(add_88_21_n_693), .b(n_2487), .y(n_2488));
nor2 g7132 (.a(n_1316), .b(n_2187), .y(n_2487));
nand2 g7134 (.a(add_88_21_n_746), .b(n_2489), .y(n_2490));
nor2 g7135 (.a(n_2846), .b(n_2189), .y(n_2489));
nand2 g53 (.a(n_1776), .b(n_2497), .y(n_2498));
nand2 g54 (.a(n_2496), .b(n_1769), .y(n_2497));
nand2 g7136 (.a(n_2495), .b(n_1758), .y(n_2496));
inv g7137 (.a(n_2494), .y(n_2495));
nand2 g7138 (.a(add_88_21_n_744), .b(add_88_21_n_787), .y(n_2494));
nand2 g7139 (.a(n_1758), .b(add_88_21_n_744), .y(n_2499));
nand2 g94 (.a(n_2500), .b(n_2505), .y(n_2506));
inv g7140 (.a(n_1797), .y(n_2500));
nand2 g7141 (.a(n_2503), .b(n_2504), .y(n_2505));
nand2 g96 (.a(n_2502), .b(n_1779), .y(n_2503));
nor2 g7142 (.a(add_88_21_n_742), .b(add_88_21_n_797), .y(n_2502));
inv g7143 (.a(n_1789), .y(n_2504));
nand2 g7144 (.a(n_1779), .b(n_3294), .y(n_2507));
nand2 g487 (.a(n_2516), .b(n_2519), .y(n_2520));
nor2 g7145 (.a(n_2513), .b(n_2515), .y(n_2516));
nor2 g7146 (.a(n_2509), .b(n_2512), .y(n_2513));
nand2 g7147 (.a(n_3936), .b(n_3953), .y(n_2509));
nand2 g7149 (.a(n_2510), .b(n_2511), .y(n_2512));
inv g7150 (.a(n_3951), .y(n_2510));
inv g7151 (.a(n_3713), .y(n_2511));
nor2 g7152 (.a(n_3952), .b(n_2511), .y(n_2515));
nor2 g7154 (.a(n_2517), .b(n_2518), .y(n_2519));
inv g7155 (.a(n_3687), .y(n_2517));
nor2 g7156 (.a(n_3936), .b(n_2511), .y(n_2518));
inv g7160 (.a(add_76_21_n_820), .y(n_2523));
inv g7163 (.a(add_76_21_n_1004), .y(n_2526));
nor2 g7167 (.a(add_76_82_n_896), .b(add_76_82_n_1092), .y(n_2531));
nand2 g7170 (.a(n_2362), .b(n_2535), .y(n_2536));
inv g7171 (.a(n_2534), .y(n_2535));
nand2 g7172 (.a(n_2579), .b(add_76_82_n_1093), .y(n_2534));
nand2 g7175 (.a(n_2546), .b(n_2551), .y(n_2552));
nor2 g7176 (.a(n_2542), .b(n_2545), .y(n_2546));
nor2 g7177 (.a(n_3843), .b(n_2541), .y(n_2542));
nand2 g424 (.a(n_1574), .b(add_76_69_n_749), .y(n_2541));
mux2 g7178 (.a(n_2544), .b(n_2543), .sel(n_1574), .y(n_2545));
nor2 g425 (.a(n_2543), .b(add_76_69_n_875), .y(n_2544));
inv g427 (.a(add_76_69_n_749), .y(n_2543));
nor2 g7179 (.a(n_2549), .b(n_2550), .y(n_2551));
nor2 g422 (.a(n_2566), .b(n_2548), .y(n_2549));
nand2 g426 (.a(n_2547), .b(add_76_69_n_875), .y(n_2548));
inv g428 (.a(n_1574), .y(n_2547));
nor2 g7180 (.a(n_2565), .b(n_2548), .y(n_2550));
nand2 g7181 (.a(n_2557), .b(n_2562), .y(n_2563));
nand2 g352 (.a(n_2554), .b(n_2556), .y(n_2557));
nor2 g360 (.a(n_2553), .b(v0_19_), .y(n_2554));
inv g361 (.a(n_2552), .y(n_2553));
nand2 g356 (.a(n_2555), .b(n_2237), .y(n_2556));
nor2 g357 (.a(n_2232), .b(n_2233), .y(n_2555));
nand2 g353 (.a(n_2558), .b(n_2561), .y(n_2562));
nor2 g359 (.a(n_2552), .b(n_2232), .y(n_2558));
inv g354 (.a(n_2560), .y(n_2561));
nand2 g355 (.a(n_2237), .b(n_2559), .y(n_2560));
nor2 g358 (.a(n_2233), .b(v0_19_), .y(n_2559));
xor2 g7182 (.a(n_2556), .b(n_2552), .y(n_2564));
xor2 g7183 (.a(n_3843), .b(n_2568), .y(n_2569));
nand2 g62 (.a(add_76_69_n_706), .b(add_76_69_n_786), .y(n_2565));
nor2 g63 (.a(add_76_69_n_729), .b(add_76_69_n_766), .y(n_2566));
xor2 g7185 (.a(add_76_82_n_1168), .b(add_76_69_n_964), .y(n_2568));
nand2 g7186 (.a(n_2571), .b(n_2575), .y(n_2576));
inv g81 (.a(n_2570), .y(n_2571));
nand2 g82 (.a(n_2807), .b(add_76_82_n_1085), .y(n_2570));
nor2 g80 (.a(n_2572), .b(n_2574), .y(n_2575));
nand2 g84 (.a(add_76_82_n_1095), .b(add_76_82_n_1084), .y(n_2572));
nand2 g86 (.a(add_76_82_n_1091), .b(n_2573), .y(n_2574));
inv g87 (.a(add_76_82_n_1232), .y(n_2573));
nor2 g77 (.a(n_2580), .b(add_76_82_n_1232), .y(n_2581));
inv g78 (.a(n_2579), .y(n_2580));
nor2 g79 (.a(n_2577), .b(n_2578), .y(n_2579));
nand2 g85 (.a(add_76_82_n_1085), .b(add_76_82_n_1095), .y(n_2577));
nand2 g83 (.a(add_76_82_n_1084), .b(add_76_82_n_1091), .y(n_2578));
mux2 g368 (.a(n_2583), .b(n_2584), .sel(n_2586), .y(n_2587));
nor2 g7187 (.a(n_2582), .b(n_1224), .y(n_2583));
inv g7188 (.a(n_2195), .y(n_2582));
nor2 g372 (.a(n_1224), .b(n_2195), .y(n_2584));
nand2 g370 (.a(n_2585), .b(n_1971), .y(n_2586));
nor2 g371 (.a(n_1956), .b(n_1964), .y(n_2585));
xor2 g369 (.a(n_2586), .b(n_2195), .y(n_2588));
nand2 g671 (.a(n_2595), .b(n_2600), .y(n_2601));
nand2 g674 (.a(n_2592), .b(n_2594), .y(n_2595));
nor2 g677 (.a(n_2589), .b(n_2591), .y(n_2592));
nand2 g682 (.a(add_76_69_n_741), .b(n_1465), .y(n_2589));
nand2 g683 (.a(add_76_69_n_759), .b(n_2590), .y(n_2591));
inv g684 (.a(v0_15_), .y(n_2590));
inv g678 (.a(n_2593), .y(n_2594));
nor2 g679 (.a(add_76_69_n_705), .b(add_76_69_n_825), .y(n_2593));
nand2 g673 (.a(n_2598), .b(n_2599), .y(n_2600));
inv g675 (.a(n_2597), .y(n_2598));
nor2 g676 (.a(n_2596), .b(n_2593), .y(n_2597));
nand2 g680 (.a(add_76_69_n_741), .b(add_76_69_n_759), .y(n_2596));
nor2 g681 (.a(n_1465), .b(v0_15_), .y(n_2599));
xor2 g672 (.a(n_2597), .b(n_1465), .y(n_2602));
xor2 g7195 (.a(n_3505), .b(n_3580), .y(n_2610));
nand2 g7197 (.a(n_2614), .b(n_2617), .y(n_2618));
nor2 g7198 (.a(n_2612), .b(add_76_82_n_898), .y(n_2614));
nor2 g7199 (.a(add_76_82_n_896), .b(add_76_82_n_980), .y(n_2612));
nand2 g7202 (.a(n_2362), .b(n_2616), .y(n_2617));
inv g7203 (.a(n_2615), .y(n_2616));
nand2 g7204 (.a(add_76_82_n_979), .b(n_2579), .y(n_2615));
nand2 g7206 (.a(n_2362), .b(n_2579), .y(n_2619));
nand2 g541 (.a(n_2625), .b(n_2629), .y(n_2630));
nand2 g544 (.a(n_2651), .b(n_2624), .y(n_2625));
nor2 g550 (.a(n_1608), .b(v0_25_), .y(n_2624));
nand2 g542 (.a(n_2633), .b(n_2628), .y(n_2629));
nor2 g545 (.a(n_2634), .b(n_2627), .y(n_2628));
nand2 g547 (.a(n_1608), .b(n_2626), .y(n_2627));
nor2 g548 (.a(add_76_69_n_1027), .b(v0_25_), .y(n_2626));
nand2 g7207 (.a(n_2638), .b(n_2648), .y(n_2649));
nand2 g7208 (.a(n_2633), .b(n_2637), .y(n_2638));
nand2 g794 (.a(n_3843), .b(add_76_69_n_753), .y(n_2633));
nor2 g796 (.a(n_2634), .b(n_2636), .y(n_2637));
nor2 g801 (.a(n_2320), .b(add_76_69_n_1043), .y(n_2634));
nand2 g803 (.a(n_1608), .b(add_76_69_n_1060), .y(n_2636));
nor2 g789 (.a(n_2642), .b(n_2647), .y(n_2648));
nor2 g795 (.a(add_76_69_n_664), .b(n_2641), .y(n_2642));
nand2 g802 (.a(n_2640), .b(add_76_69_n_753), .y(n_2641));
inv g805 (.a(n_1608), .y(n_2640));
nand2 g7209 (.a(n_2645), .b(n_2646), .y(n_2647));
nand2 g797 (.a(n_2321), .b(n_2644), .y(n_2645));
nor2 g800 (.a(n_1608), .b(add_76_69_n_1043), .y(n_2644));
nand2 g804 (.a(n_2640), .b(add_76_69_n_1027), .y(n_2646));
nand2 g7210 (.a(n_2633), .b(n_2650), .y(n_2651));
nor2 g793 (.a(n_2634), .b(add_76_69_n_1027), .y(n_2650));
nand2 g145 (.a(n_2654), .b(n_2656), .y(n_2657));
inv g7211 (.a(n_2653), .y(n_2654));
nor2 g7212 (.a(n_2652), .b(add_76_82_n_1299), .y(n_2653));
nor2 g148 (.a(add_76_82_n_915), .b(add_76_82_n_959), .y(n_2652));
nor2 g149 (.a(add_76_82_n_1211), .b(v0_25_), .y(n_2656));
nor2 g144 (.a(n_2653), .b(add_76_82_n_1211), .y(n_2658));
nand2 g7215 (.a(n_2660), .b(n_2662), .y(n_2663));
nor2 g7216 (.a(n_2659), .b(v0_27_), .y(n_2660));
inv g7217 (.a(n_1668), .y(n_2659));
nand2 g7218 (.a(n_2661), .b(add_76_82_n_864), .y(n_2662));
nand2 g7219 (.a(n_3866), .b(add_76_82_n_963), .y(n_2661));
nand2 g7220 (.a(n_2666), .b(n_2661), .y(n_2667));
nor2 g7221 (.a(n_1668), .b(n_2665), .y(n_2666));
nand2 g7222 (.a(add_76_82_n_864), .b(n_2664), .y(n_2665));
inv g7223 (.a(v0_27_), .y(n_2664));
xor2 g7224 (.a(n_2662), .b(n_1668), .y(n_2669));
nor2 g7225 (.a(n_2671), .b(n_2674), .y(n_2675));
nand2 g7226 (.a(n_2670), .b(add_76_21_n_891), .y(n_2671));
inv g7227 (.a(add_76_21_n_811), .y(n_2670));
nor2 g7228 (.a(n_3941), .b(n_2673), .y(n_2674));
inv g7230 (.a(add_76_21_n_948), .y(n_2673));
nor2 g45 (.a(n_2903), .b(n_2682), .y(n_2683));
inv g7232 (.a(n_2681), .y(n_2682));
nor2 g47 (.a(n_2680), .b(sum_2_), .y(n_2681));
inv g48 (.a(n_2679), .y(n_2680));
nor2 g49 (.a(n_496), .b(n_494), .y(n_2679));
nand2 g7233 (.a(n_2688), .b(n_2692), .y(n_2693));
nand2 g7234 (.a(n_2873), .b(n_2687), .y(n_2688));
nand2 g7237 (.a(n_2686), .b(add_76_82_n_1210), .y(n_2687));
nand2 g7238 (.a(n_1846), .b(n_1850), .y(n_2686));
nand2 g7239 (.a(n_2877), .b(n_2686), .y(n_2692));
nand2 g7241 (.a(add_76_82_n_1210), .b(n_2689), .y(n_2690));
inv g7242 (.a(v0_5_), .y(n_2689));
inv g7244 (.a(n_3913), .y(n_2696));
nor2 g7248 (.a(n_2911), .b(n_2704), .y(n_2705));
nor2 g7249 (.a(n_2792), .b(n_2793), .y(n_2704));
inv g289 (.a(add_76_82_n_1144), .y(n_2702));
nand2 g7252 (.a(n_2712), .b(n_2716), .y(n_2717));
nand2 g7253 (.a(n_2709), .b(n_2711), .y(n_2712));
nor2 g7254 (.a(n_2708), .b(v0_7_), .y(n_2709));
inv g7255 (.a(n_1517), .y(n_2708));
nand2 g7256 (.a(n_3910), .b(add_76_82_n_960), .y(n_2711));
nand2 g7258 (.a(n_2715), .b(n_3910), .y(n_2716));
nor2 g7259 (.a(n_1517), .b(n_2714), .y(n_2715));
nand2 g7260 (.a(add_76_82_n_960), .b(n_2713), .y(n_2714));
inv g7261 (.a(v0_7_), .y(n_2713));
xor2 g7262 (.a(n_2711), .b(n_1517), .y(n_2718));
nand2 g7263 (.a(n_2724), .b(n_2729), .y(n_2730));
nand2 g7264 (.a(n_2720), .b(n_4048), .y(n_2724));
nor2 g7265 (.a(n_3580), .b(n_2719), .y(n_2720));
inv g7266 (.a(n_3272), .y(n_2719));
nand2 g7270 (.a(n_2726), .b(n_2728), .y(n_2729));
nor2 g7271 (.a(n_3580), .b(n_2725), .y(n_2726));
nand2 g7272 (.a(n_1890), .b(n_2719), .y(n_2725));
nor2 g7273 (.a(n_4049), .b(n_3668), .y(n_2728));
xor2 g7275 (.a(n_4048), .b(n_3272), .y(n_2731));
nand2 g7276 (.a(n_2736), .b(n_2740), .y(n_2741));
nand2 g7277 (.a(n_2734), .b(n_2735), .y(n_2736));
inv g7278 (.a(n_2733), .y(n_2734));
nor2 g7279 (.a(n_2732), .b(add_76_69_n_755), .y(n_2733));
nor2 g7280 (.a(add_76_69_n_705), .b(add_76_69_n_872), .y(n_2732));
nor2 g7281 (.a(n_1490), .b(v0_11_), .y(n_2735));
inv g7282 (.a(n_2739), .y(n_2740));
nor2 g7283 (.a(n_2738), .b(n_2732), .y(n_2739));
nand2 g7284 (.a(n_2737), .b(n_1490), .y(n_2738));
nor2 g7285 (.a(add_76_69_n_755), .b(v0_11_), .y(n_2737));
inv g7289 (.a(add_76_21_n_859), .y(n_2743));
nand2 g7294 (.a(n_2749), .b(add_76_21_n_1038), .y(n_2750));
inv g7295 (.a(add_76_21_n_815), .y(n_2749));
nor2 g7296 (.a(n_3941), .b(add_76_21_n_1071), .y(n_2753));
nor2 g30 (.a(n_2060), .b(n_2755), .y(n_2756));
inv g33 (.a(sum_0_), .y(n_2755));
nor2 g7299 (.a(n_2755), .b(sum_1_), .y(n_2757));
nor2 g7300 (.a(n_2755), .b(n_179), .y(n_2758));
nand2 g1150 (.a(n_2251), .b(n_2760), .y(n_2761));
nor2 g1155 (.a(n_2759), .b(v0_17_), .y(n_2760));
inv g1156 (.a(n_2256), .y(n_2759));
nor2 g1148 (.a(n_2764), .b(n_2765), .y(n_2766));
nand2 g1153 (.a(n_2762), .b(n_2763), .y(n_2764));
inv g1158 (.a(n_2262), .y(n_2762));
inv g1157 (.a(n_3908), .y(n_2763));
nor2 g1154 (.a(add_76_82_n_896), .b(add_76_82_n_1232), .y(n_2765));
nor2 g1145 (.a(n_2770), .b(n_2765), .y(n_2771));
nand2 g1149 (.a(n_2762), .b(n_2769), .y(n_2770));
nor2 g1152 (.a(n_3908), .b(v0_17_), .y(n_2769));
nand2 g1151 (.a(n_2251), .b(n_2256), .y(n_2772));
inv g7312 (.a(n_4350), .y(n_2792));
nand2 g7313 (.a(n_2702), .b(n_2915), .y(n_2793));
nand2 g195 (.a(add_76_82_n_1081), .b(add_76_82_n_1088), .y(n_2798));
nor2 g188 (.a(n_2798), .b(add_76_82_n_1208), .y(n_2805));
inv g194 (.a(n_2798), .y(n_2807));
nand2 g668 (.a(n_2813), .b(n_2814), .y(n_2815));
nand2 g7315 (.a(add_76_21_n_902), .b(n_2812), .y(n_2813));
inv g7316 (.a(n_1827), .y(n_2812));
nand2 g7317 (.a(n_2812), .b(add_76_21_n_1249), .y(n_2814));
inv g659 (.a(n_2820), .y(n_2821));
nand2 g660 (.a(n_2816), .b(n_2819), .y(n_2820));
nor2 g7318 (.a(add_76_21_n_902), .b(n_3709), .y(n_2816));
nor2 g667 (.a(n_3664), .b(n_2818), .y(n_2819));
inv g7319 (.a(n_2817), .y(n_2818));
nor2 g7320 (.a(n_2812), .b(add_76_21_n_1249), .y(n_2817));
nor2 g662 (.a(n_3710), .b(n_2824), .y(n_2825));
nand2 g664 (.a(n_2823), .b(n_2812), .y(n_2824));
nor2 g670 (.a(add_76_21_n_1011), .b(n_1551), .y(n_2823));
nor2 g661 (.a(add_76_21_n_902), .b(n_2827), .y(n_2828));
nand2 g663 (.a(n_2826), .b(n_2817), .y(n_2827));
inv g669 (.a(n_2823), .y(n_2826));
nand2 g665 (.a(add_76_21_n_942), .b(n_2831), .y(n_2832));
inv g7321 (.a(n_3710), .y(n_2831));
nand2 g666 (.a(n_2831), .b(add_76_21_n_949), .y(n_2833));
inv g7324 (.a(n_4088), .y(n_2841));
nor2 g7329 (.a(n_2587), .b(n_4088), .y(n_2842));
nor2 g7330 (.a(n_3956), .b(n_4088), .y(n_2843));
nor2 g7333 (.a(add_88_21_n_865), .b(add_88_21_n_882), .y(n_2846));
nand2 g7339 (.a(add_88_21_n_747), .b(n_3892), .y(n_2852));
nor2 g7340 (.a(n_2125), .b(n_4031), .y(n_2853));
inv g7341 (.a(n_4031), .y(n_2854));
nor2 g423 (.a(n_2868), .b(n_2690), .y(n_2862));
mux2 g474 (.a(n_2867), .b(n_2869), .sel(n_2872), .y(n_2873));
nor2 g478 (.a(n_2866), .b(v0_5_), .y(n_2867));
nand2 g482 (.a(add_76_69_n_734), .b(add_76_69_n_1021), .y(n_2866));
nor2 g480 (.a(n_2868), .b(v0_5_), .y(n_2869));
inv g481 (.a(n_2866), .y(n_2868));
xor2 g477 (.a(n_2870), .b(n_2871), .y(n_2872));
nor2 g484 (.a(add_76_82_n_1257), .b(add_76_82_n_1273), .y(n_2870));
nor2 g483 (.a(add_76_69_n_997), .b(add_76_69_n_1078), .y(n_2871));
xor2 g473 (.a(n_2687), .b(n_2874), .y(n_2875));
xor2 g476 (.a(n_2872), .b(n_2866), .y(n_2874));
mux2 g475 (.a(n_2862), .b(n_2876), .sel(n_2872), .y(n_2877));
nor2 g479 (.a(n_2866), .b(n_2690), .y(n_2876));
inv g107 (.a(n_2880), .y(n_2881));
nor2 g108 (.a(n_2878), .b(n_2879), .y(n_2880));
nand2 g110 (.a(n_395), .b(n_281), .y(n_2878));
nand2 g7353 (.a(n_344), .b(n_379), .y(n_2879));
nand2 g7363 (.a(n_2680), .b(sum_2_), .y(n_2901));
nand2 g347 (.a(n_2902), .b(n_2901), .y(n_2903));
nand2 g7366 (.a(n_2881), .b(sum_3_), .y(n_2902));
inv g7367 (.a(n_2904), .y(n_2905));
nor2 g7368 (.a(n_2881), .b(sum_3_), .y(n_2904));
inv g7370 (.a(n_2910), .y(n_2911));
nand2 g7371 (.a(n_2909), .b(n_2903), .y(n_2910));
nor2 g350 (.a(add_76_82_n_1144), .b(n_2904), .y(n_2909));
inv g7372 (.a(n_2902), .y(n_2912));
nand2 g348 (.a(n_1870), .b(n_2902), .y(n_2914));
nor2 g7373 (.a(n_2681), .b(n_2904), .y(n_2915));
nor2 g7374 (.a(n_2693), .b(n_2921), .y(n_2922));
mux2 g7375 (.a(n_2918), .b(n_2919), .sel(n_2920), .y(n_2921));
nand2 g7376 (.a(n_2917), .b(v0_4_), .y(n_2918));
inv g7377 (.a(n_2916), .y(n_2917));
xor2 g236 (.a(n_2927), .b(add_76_69_n_995), .y(n_2916));
nand2 g7378 (.a(n_2916), .b(v0_4_), .y(n_2919));
nand2 g237 (.a(n_3912), .b(n_2705), .y(n_2920));
inv g7379 (.a(n_2921), .y(n_2923));
nand2 g228 (.a(add_76_21_n_889), .b(n_2921), .y(n_2924));
nor2 g7380 (.a(n_2925), .b(v0_4_), .y(n_2926));
xor2 g7381 (.a(n_2920), .b(n_2916), .y(n_2925));
nand2 g7382 (.a(add_76_69_n_815), .b(add_76_69_n_874), .y(n_2927));
nand2 g745 (.a(n_2933), .b(n_2940), .y(n_2941));
nand2 g7383 (.a(n_2929), .b(n_2932), .y(n_2933));
nand2 g7384 (.a(n_2927), .b(n_2928), .y(n_2929));
nor2 g760 (.a(add_76_69_n_1078), .b(add_76_69_n_1023), .y(n_2928));
nor2 g754 (.a(n_2931), .b(add_76_69_n_913), .y(n_2932));
nand2 g7385 (.a(add_76_69_n_977), .b(add_76_69_n_1044), .y(n_2931));
nor2 g746 (.a(n_2935), .b(n_2939), .y(n_2940));
nor2 g749 (.a(n_2934), .b(add_76_69_n_977), .y(n_2935));
nor2 g756 (.a(add_76_69_n_913), .b(add_76_69_n_997), .y(n_2934));
nor2 g7387 (.a(add_76_69_n_748), .b(n_2938), .y(n_2939));
nand2 g7389 (.a(n_2937), .b(n_2928), .y(n_2938));
inv g7390 (.a(add_76_69_n_977), .y(n_2937));
inv g7391 (.a(n_2934), .y(n_2942));
nor2 g751 (.a(n_2934), .b(add_76_69_n_1101), .y(n_2943));
nand2 g7392 (.a(add_76_69_n_890), .b(n_2928), .y(n_2944));
inv g759 (.a(n_2928), .y(n_2945));
nor2 g7393 (.a(add_76_21_n_881), .b(add_76_21_n_930), .y(n_2946));
nand2 g729 (.a(n_2953), .b(n_2960), .y(n_2961));
nand2 g731 (.a(n_2949), .b(n_2952), .y(n_2953));
nand2 g738 (.a(n_2947), .b(n_3699), .y(n_2949));
inv g7394 (.a(n_2946), .y(n_2947));
nor2 g7396 (.a(n_2950), .b(n_3677), .y(n_2952));
nand2 g7397 (.a(add_76_21_n_1144), .b(n_2019), .y(n_2950));
nor2 g730 (.a(n_2956), .b(n_2959), .y(n_2960));
nor2 g732 (.a(n_2946), .b(n_2955), .y(n_2956));
nand2 g7399 (.a(n_2954), .b(n_3699), .y(n_2955));
inv g7400 (.a(add_76_21_n_1144), .y(n_2954));
nor2 g736 (.a(n_2958), .b(add_76_21_n_1144), .y(n_2959));
inv g7401 (.a(n_3679), .y(n_2958));
nand2 g7403 (.a(add_76_21_n_957), .b(n_2947), .y(n_2963));
nand2 g735 (.a(n_3699), .b(n_4399), .y(n_2966));
xor2 add_88_82_g7421 (.a(v1_31_), .b(n_2981), .y(n_2982));
xor2 add_88_82_g7422 (.a(n_687), .b(n_1280), .y(n_2981));
nand2 add_88_82_g7423 (.a(add_88_82_n_1889), .b(add_88_82_n_2196), .y(n_2983));
nand2 add_88_82_g7431 (.a(add_88_82_n_1893), .b(add_88_82_n_2188), .y(n_2993));
xor2 g6430__7432 (.a(n_2997), .b(n_1459), .y(n_2998));
xor2 add_88_69_g1531__7433 (.a(n_2996), .b(n_2993), .y(n_2997));
xor2 add_88_82_g7434 (.a(n_2994), .b(n_2995), .y(n_2996));
nor2 add_88_69_g7435 (.a(add_88_69_n_1697), .b(add_88_69_n_1649), .y(n_2994));
xor2 add_88_82_g7436 (.a(n_686), .b(n_1281), .y(n_2995));
nor2 g7443 (.a(n_3983), .b(v0_28_), .y(n_3010));
nand2 add_76_82_g7448 (.a(add_76_82_n_850), .b(add_76_82_n_856), .y(n_3008));
nand2 g7449 (.a(n_3983), .b(v0_28_), .y(n_3011));
nor2 g7534 (.a(n_653), .b(n_3110), .y(n_3111));
nand2 g7536 (.a(n_181), .b(n_3109), .y(n_3110));
inv g7537 (.a(counter_3_), .y(n_3109));
nand2 g7538 (.a(n_192), .b(n_181), .y(n_3112));
nand2 g7549 (.a(n_688), .b(sum_0_), .y(n_3125));
nor2 add_76_21_g7550 (.a(n_3129), .b(v0_1_), .y(n_3130));
xor2 g6397__7551 (.a(n_3127), .b(n_3128), .y(n_3129));
xor2 add_76_82_g7552 (.a(n_3126), .b(n_3125), .y(n_3127));
xor2 add_76_69_g7553 (.a(add_76_69_n_983), .b(add_76_69_n_1013), .y(n_3126));
nand2 add_76_82_g7554 (.a(n_1861), .b(add_76_82_n_1196), .y(n_3128));
nand2 add_76_21_g7555 (.a(n_3129), .b(v0_1_), .y(n_3131));
nand2 g35 (.a(add_76_21_n_951), .b(n_2947), .y(n_3134));
xor2 add_76_21_g7558 (.a(n_2924), .b(add_76_21_n_1158), .y(n_3139));
xor2 add_88_21_g7560 (.a(n_3143), .b(v1_0_), .y(n_3144));
xor2 g6442__7561 (.a(n_3142), .b(n_3139), .y(n_3143));
xor2 add_88_69_g7562 (.a(n_3141), .b(n_3269), .y(n_3142));
nor2 add_88_82_g7563 (.a(n_2062), .b(n_2756), .y(n_3141));
nand2 add_88_21_g7564 (.a(n_3143), .b(v1_0_), .y(n_3145));
nand2 add_88_69_g7576 (.a(n_3139), .b(n_3269), .y(n_3157));
nor2 add_88_21_g7577 (.a(n_3161), .b(v1_1_), .y(n_3162));
xor2 g6441__7578 (.a(n_3159), .b(n_3160), .y(n_3161));
xor2 add_88_69_g1713__7579 (.a(n_3158), .b(n_3157), .y(n_3159));
xor2 add_88_82_g7580 (.a(add_88_82_n_2139), .b(n_2062), .y(n_3158));
nand2 add_88_69_g7581 (.a(add_88_69_n_1703), .b(add_88_69_n_1635), .y(n_3160));
nand2 add_88_21_g7582 (.a(n_3161), .b(v1_1_), .y(n_3163));
nand2 add_88_69_g1752__7583 (.a(add_88_69_n_1514), .b(add_88_69_n_1703), .y(n_3164));
nor2 add_88_21_g7584 (.a(n_3168), .b(v1_2_), .y(n_3169));
xor2 g6444__7585 (.a(n_3167), .b(n_3164), .y(n_3168));
xor2 add_88_69_g1671__7586 (.a(n_3165), .b(n_3166), .y(n_3167));
nor2 add_88_69_g7587 (.a(add_88_69_n_1645), .b(add_88_69_n_1729), .y(n_3165));
xor2 add_88_82_g7588 (.a(n_2078), .b(add_88_82_n_2138), .y(n_3166));
nand2 add_88_21_g7589 (.a(n_3168), .b(v1_2_), .y(n_3170));
nor2 g7593 (.a(add_88_21_n_1014), .b(n_4371), .y(n_3172));
nand2 g7597 (.a(n_4371), .b(v1_r_6_), .y(n_3177));
nor2 add_88_21_g7598 (.a(n_3183), .b(v1_3_), .y(n_3184));
xor2 g6395__7599 (.a(n_3181), .b(n_3182), .y(n_3183));
xor2 add_88_69_g1628__7600 (.a(n_3179), .b(n_3180), .y(n_3181));
xor2 add_88_82_g7601 (.a(add_88_82_n_2010), .b(add_88_82_n_2137), .y(n_3179));
nor2 add_88_69_g7602 (.a(add_88_69_n_1698), .b(add_88_69_n_1718), .y(n_3180));
nand2 add_88_69_g1678__7603 (.a(add_88_69_n_1452), .b(add_88_69_n_1644), .y(n_3182));
nand2 add_88_21_g7604 (.a(n_3183), .b(v1_3_), .y(n_3185));
nor2 add_88_21_g7605 (.a(n_3190), .b(v1_5_), .y(n_3191));
xor2 g6393__7606 (.a(n_3188), .b(n_3189), .y(n_3190));
xor2 add_88_69_g1605__7607 (.a(n_3186), .b(n_3187), .y(n_3188));
xor2 add_88_82_g7608 (.a(add_88_82_n_1994), .b(add_88_82_n_2136), .y(n_3186));
nor2 add_88_69_g7609 (.a(add_88_69_n_1700), .b(add_88_69_n_1646), .y(n_3187));
nand2 add_88_69_g1634__7610 (.a(add_88_69_n_1355), .b(add_88_69_n_1728), .y(n_3189));
nand2 add_88_21_g7611 (.a(n_3190), .b(v1_5_), .y(n_3192));
nor2 g7615 (.a(add_88_21_n_1008), .b(n_4371), .y(n_3194));
nand2 g7619 (.a(n_4371), .b(v1_r_10_), .y(n_3199));
xor2 add_88_69_g1588__7622 (.a(n_3201), .b(n_3202), .y(n_3203));
xor2 add_88_82_g7623 (.a(add_88_82_n_1981), .b(add_88_82_n_2134), .y(n_3201));
nor2 add_88_69_g7624 (.a(add_88_69_n_1711), .b(add_88_69_n_1653), .y(n_3202));
nand2 add_88_69_g1609__7625 (.a(add_88_69_n_1397), .b(add_88_69_n_1323), .y(n_3204));
nand2 add_88_21_g7626 (.a(n_3337), .b(v1_7_), .y(n_3207));
nor2 g7630 (.a(add_88_21_n_992), .b(n_4371), .y(n_3209));
nand2 g7634 (.a(n_4371), .b(v1_r_9_), .y(n_3214));
nor2 g7638 (.a(add_88_21_n_1010), .b(n_4371), .y(n_3217));
nand2 g7642 (.a(n_4371), .b(v1_r_12_), .y(n_3222));
nor2 g7646 (.a(add_88_21_n_1015), .b(n_4371), .y(n_3225));
nand2 g7650 (.a(n_4371), .b(v1_r_11_), .y(n_3230));
nor2 g7651 (.a(n_3232), .b(add_88_21_n_758), .y(n_3233));
nand2 g7652 (.a(n_2179), .b(n_3284), .y(n_3232));
nor2 g38 (.a(n_3434), .b(n_3236), .y(n_3237));
inv g40 (.a(add_88_21_n_896), .y(n_3236));
nor2 g7657 (.a(add_88_21_n_999), .b(n_4371), .y(n_3239));
nand2 g7661 (.a(n_4371), .b(v1_r_15_), .y(n_3244));
nor2 g7665 (.a(add_88_21_n_979), .b(n_4371), .y(n_3247));
nand2 g7669 (.a(n_4371), .b(v1_r_14_), .y(n_3252));
nor2 g7673 (.a(add_88_21_n_1000), .b(n_4371), .y(n_3255));
nand2 g7677 (.a(n_4371), .b(v1_r_13_), .y(n_3260));
xor2 add_76_82_g7680 (.a(n_3262), .b(n_3263), .y(n_3264));
xor2 add_76_69_g7681 (.a(add_76_69_n_778), .b(add_76_69_n_954), .y(n_3262));
nor2 g7682 (.a(n_2912), .b(n_2904), .y(n_3263));
nand2 add_76_82_g7683 (.a(n_1868), .b(n_2901), .y(n_3265));
nand2 add_76_21_g7684 (.a(n_3319), .b(v0_3_), .y(n_3268));
xor2 g71 (.a(add_76_21_n_837), .b(n_3270), .y(n_3271));
xor2 g7685 (.a(add_76_21_n_1141), .b(n_3269), .y(n_3270));
xor2 g7686 (.a(n_848), .b(v0_0_), .y(n_3269));
xor2 g7687 (.a(add_76_21_n_837), .b(add_76_21_n_1141), .y(n_3272));
nor2 add_88_21_g7688 (.a(n_3277), .b(v1_9_), .y(n_3278));
xor2 g6392__7689 (.a(n_3275), .b(n_3276), .y(n_3277));
xor2 add_88_69_g1552__7690 (.a(n_3273), .b(n_3274), .y(n_3275));
xor2 add_88_82_g7691 (.a(add_88_82_n_1952), .b(add_88_82_n_2132), .y(n_3273));
nor2 add_88_69_g7692 (.a(add_88_69_n_1701), .b(add_88_69_n_1714), .y(n_3274));
nand2 add_88_69_g1582__7693 (.a(add_88_69_n_1288), .b(add_88_69_n_1723), .y(n_3276));
nand2 add_88_21_g7694 (.a(n_3277), .b(v1_9_), .y(n_3279));
nor2 g7698 (.a(n_3283), .b(add_88_21_n_805), .y(n_3284));
nor2 g7699 (.a(n_3434), .b(add_88_21_n_887), .y(n_3283));
mux2 g7704 (.a(n_3290), .b(n_3291), .sel(n_1541), .y(n_3292));
nor2 g7705 (.a(n_3289), .b(v1_19_), .y(n_3290));
inv g7706 (.a(n_1540), .y(n_3289));
nor2 g7707 (.a(n_1540), .b(v1_19_), .y(n_3291));
xor2 g7708 (.a(n_1541), .b(n_1540), .y(n_3293));
inv fopt7709 (.a(add_88_21_n_742), .y(n_3294));
mux2 g7710 (.a(n_3297), .b(n_3298), .sel(n_1484), .y(n_3299));
nor2 g7711 (.a(n_3296), .b(v1_21_), .y(n_3297));
inv g7712 (.a(n_1483), .y(n_3296));
nor2 g7713 (.a(n_1483), .b(v1_21_), .y(n_3298));
xor2 g7714 (.a(n_1484), .b(n_1483), .y(n_3300));
nand2 g7726 (.a(n_3134), .b(n_1414), .y(n_3311));
mux2 g7729 (.a(n_3316), .b(n_3317), .sel(n_3264), .y(n_3318));
nor2 g7730 (.a(n_3315), .b(v0_3_), .y(n_3316));
inv g7731 (.a(n_3265), .y(n_3315));
nor2 g7732 (.a(n_3265), .b(v0_3_), .y(n_3317));
xor2 g7733 (.a(n_3264), .b(n_3265), .y(n_3319));
nor2 add_88_21_g7734 (.a(n_3324), .b(v1_6_), .y(n_3325));
xor2 g6440__7735 (.a(n_3322), .b(n_3323), .y(n_3324));
xor2 add_88_69_g1604__7736 (.a(n_3320), .b(n_3321), .y(n_3322));
xor2 add_88_82_g7737 (.a(add_88_82_n_1989), .b(add_88_82_n_2135), .y(n_3320));
nor2 add_88_69_g7738 (.a(add_88_69_n_1654), .b(add_88_69_n_1674), .y(n_3321));
nand2 add_88_69_g1635__7739 (.a(add_88_69_n_1501), .b(add_88_69_n_1342), .y(n_3323));
nand2 add_88_21_g7740 (.a(n_3324), .b(v1_6_), .y(n_3326));
mux2 g7741 (.a(n_3328), .b(n_3330), .sel(n_3331), .y(n_3332));
nand2 g7612_dup2 (.a(n_3327), .b(n_3199), .y(n_3328));
inv g7742 (.a(n_3194), .y(n_3327));
nand2 g7743 (.a(n_3329), .b(n_3199), .y(n_3330));
nand2 g7744 (.a(add_88_21_n_1008), .b(n_1683), .y(n_3329));
nand2 add_88_21_g7745 (.a(add_88_21_n_718), .b(add_88_21_n_877), .y(n_3331));
mux2 g7746 (.a(n_3334), .b(n_3335), .sel(n_3204), .y(n_3336));
nor2 g7747 (.a(n_3333), .b(v1_7_), .y(n_3334));
inv g7748 (.a(n_3203), .y(n_3333));
nor2 g7749 (.a(n_3203), .b(v1_7_), .y(n_3335));
xor2 g7750 (.a(n_3204), .b(n_3203), .y(n_3337));
mux2 g7751 (.a(n_3339), .b(n_3341), .sel(n_3342), .y(n_3343));
nand2 g7627_dup2 (.a(n_3338), .b(n_3214), .y(n_3339));
inv g7752 (.a(n_3209), .y(n_3338));
nand2 g7753 (.a(n_3340), .b(n_3214), .y(n_3341));
nand2 g7754 (.a(add_88_21_n_992), .b(n_1683), .y(n_3340));
nand2 add_88_21_g7755 (.a(add_88_21_n_715), .b(add_88_21_n_1113), .y(n_3342));
mux2 g7756 (.a(n_3345), .b(n_3347), .sel(n_3348), .y(n_3349));
nand2 g7643_dup2 (.a(n_3344), .b(n_3230), .y(n_3345));
inv g7757 (.a(n_3225), .y(n_3344));
nand2 g7758 (.a(n_3346), .b(n_3230), .y(n_3347));
nand2 g7759 (.a(add_88_21_n_1015), .b(n_1683), .y(n_3346));
nor2 add_88_21_g7760 (.a(add_88_21_n_800), .b(add_88_21_n_721), .y(n_3348));
mux2 g7761 (.a(n_3351), .b(n_3353), .sel(n_3434), .y(n_3355));
nand2 g7635_dup2 (.a(n_3350), .b(n_3222), .y(n_3351));
inv g7762 (.a(n_3217), .y(n_3350));
nand2 g7763 (.a(n_3352), .b(n_3222), .y(n_3353));
nand2 g7764 (.a(add_88_21_n_1010), .b(n_1683), .y(n_3352));
mux2 g7766 (.a(n_3357), .b(n_3359), .sel(n_3360), .y(n_3361));
nand2 g7662_dup2 (.a(n_3356), .b(n_3252), .y(n_3357));
inv g7767 (.a(n_3247), .y(n_3356));
nand2 g7768 (.a(n_3358), .b(n_3252), .y(n_3359));
nand2 g7769 (.a(add_88_21_n_979), .b(n_1683), .y(n_3358));
nor2 add_88_21_g7770 (.a(add_88_21_n_751), .b(add_88_21_n_720), .y(n_3360));
nor2 add_88_21_g7771 (.a(n_3366), .b(v1_11_), .y(n_3367));
xor2 g6437__7772 (.a(n_3364), .b(n_3365), .y(n_3366));
xor2 add_88_69_g1554__7773 (.a(n_3362), .b(n_3363), .y(n_3364));
xor2 add_88_82_g7774 (.a(add_88_82_n_1974), .b(add_88_82_n_2120), .y(n_3362));
nand2 add_88_69_g7775 (.a(add_88_69_n_1709), .b(add_88_69_n_1719), .y(n_3363));
nor2 add_88_69_g1586__7776 (.a(add_88_69_n_1372), .b(add_88_69_n_1304), .y(n_3365));
nand2 add_88_21_g7777 (.a(n_3366), .b(v1_11_), .y(n_3368));
nand2 g7670_dup2 (.a(n_3369), .b(n_3260), .y(n_3370));
inv g7779 (.a(n_3255), .y(n_3369));
nand2 g7780 (.a(n_3371), .b(n_3260), .y(n_3372));
nand2 g7781 (.a(add_88_21_n_1000), .b(n_1683), .y(n_3371));
mux2 g7783 (.a(n_3376), .b(n_3378), .sel(n_3379), .y(n_3380));
nand2 g7654_dup2 (.a(n_3375), .b(n_3244), .y(n_3376));
inv g7784 (.a(n_3239), .y(n_3375));
nand2 g7785 (.a(n_3377), .b(n_3244), .y(n_3378));
nand2 g7786 (.a(add_88_21_n_999), .b(n_1683), .y(n_3377));
nor2 add_88_21_g7787 (.a(n_3237), .b(add_88_21_n_788), .y(n_3379));
nor2 add_88_21_g7804 (.a(n_3403), .b(v1_13_), .y(n_3404));
xor2 g6435__7805 (.a(n_3401), .b(n_3402), .y(n_3403));
xor2 add_88_69_g1558__7806 (.a(n_3399), .b(n_3400), .y(n_3401));
xor2 add_88_82_g7807 (.a(add_88_82_n_1940), .b(add_88_82_n_2128), .y(n_3399));
nor2 add_88_69_g7808 (.a(add_88_69_n_1710), .b(n_2730), .y(n_3400));
nand2 add_88_69_g1583__7809 (.a(add_88_69_n_1331), .b(add_88_69_n_1295), .y(n_3402));
nand2 add_88_21_g7810 (.a(n_3403), .b(v1_13_), .y(n_3405));
nand2 add_88_21_g7821 (.a(n_3422), .b(v1_10_), .y(n_3423));
xor2 g6438__7822 (.a(n_3420), .b(n_3421), .y(n_3422));
xor2 add_88_69_g1553__7823 (.a(n_3418), .b(n_3419), .y(n_3420));
xor2 add_88_82_g7824 (.a(add_88_82_n_1932), .b(add_88_82_n_2116), .y(n_3418));
nor2 add_88_69_g7825 (.a(add_88_69_n_1642), .b(add_88_69_n_1672), .y(n_3419));
nand2 add_88_69_g1584__7826 (.a(add_88_69_n_1297), .b(add_88_69_n_1471), .y(n_3421));
nor2 add_88_21_g7827 (.a(n_3422), .b(v1_10_), .y(n_3424));
nor2 add_88_21_g7837 (.a(add_88_21_n_781), .b(add_88_21_n_713), .y(n_3434));
inv g7838 (.a(n_3435), .y(n_3436));
nand2 g7839 (.a(add_88_21_n_860), .b(n_2179), .y(n_3435));
nand2 g7840 (.a(n_3437), .b(add_76_21_n_949), .y(n_3438));
nor2 g7841 (.a(n_3710), .b(add_76_21_n_977), .y(n_3437));
nand2 g7842 (.a(n_3439), .b(n_2353), .y(n_3440));
nor2 g7843 (.a(add_76_82_n_1034), .b(n_3907), .y(n_3439));
nor2 g7844 (.a(n_3441), .b(n_4371), .y(n_3442));
mux2 g7845 (.a(v1_26_), .b(n_1737), .sel(n_2119), .y(n_3441));
nor2 g7846 (.a(n_3443), .b(n_1998), .y(n_3444));
xor2 g7847 (.a(n_3681), .b(n_2007), .y(n_3443));
nand2 g7854 (.a(n_3451), .b(n_2142), .y(n_3452));
nor2 g7855 (.a(n_2384), .b(n_2380), .y(n_3451));
nor2 g7856 (.a(n_3453), .b(n_3490), .y(n_3454));
xor2 g7857 (.a(n_3503), .b(n_3579), .y(n_3453));
nand2 g1140 (.a(n_3487), .b(n_3489), .y(n_3490));
nor2 g7890 (.a(n_1983), .b(n_1987), .y(n_3487));
inv g7891 (.a(n_3488), .y(n_3489));
nand2 g7892 (.a(n_1990), .b(n_1991), .y(n_3488));
nand2 g7893 (.a(n_1663), .b(add_76_21_n_1203), .y(n_3491));
nor2 g7894 (.a(n_2750), .b(n_2753), .y(n_3493));
xor2 g1137 (.a(n_3493), .b(n_3491), .y(n_3502));
xor2 g857 (.a(n_3503), .b(n_3504), .y(n_3505));
nor2 g864 (.a(add_76_21_n_817), .b(add_76_21_n_882), .y(n_3503));
nand2 g861 (.a(n_1638), .b(add_76_21_n_1272), .y(n_3504));
xor2 g856 (.a(n_4048), .b(n_3524), .y(n_3514));
xor2 g7900 (.a(n_3520), .b(n_3524), .y(n_3525));
nor2 g7901 (.a(n_3518), .b(n_3519), .y(n_3520));
nand2 g7902 (.a(n_2523), .b(add_76_21_n_922), .y(n_3518));
nor2 g351 (.a(n_3941), .b(n_2526), .y(n_3519));
nand2 g7903 (.a(n_3521), .b(n_3523), .y(n_3524));
nand2 g7904 (.a(n_2669), .b(v0_27_), .y(n_3521));
inv g7905 (.a(n_3522), .y(n_3523));
nand2 g7906 (.a(n_2663), .b(n_2667), .y(n_3522));
nand2 g7909 (.a(n_3710), .b(n_1882), .y(n_3527));
nor2 g7910 (.a(n_2587), .b(n_3574), .y(n_3575));
mux2 g7911 (.a(n_3572), .b(n_3573), .sel(n_3525), .y(n_3574));
nand2 g7912 (.a(n_3505), .b(n_3571), .y(n_3572));
nand2 g7914 (.a(n_3505), .b(n_4048), .y(n_3573));
xor2 g7915 (.a(n_3577), .b(n_3578), .y(n_3579));
inv g7916 (.a(n_3576), .y(n_3577));
nor2 g313 (.a(n_3311), .b(add_76_21_n_905), .y(n_3576));
xor2 g311 (.a(n_3504), .b(add_76_21_n_1135), .y(n_3578));
xor2 g7917 (.a(n_3577), .b(add_76_21_n_1135), .y(n_3580));
inv g7922 (.a(n_3596), .y(n_3597));
nor2 g7923 (.a(n_3592), .b(n_3595), .y(n_3596));
nand2 g7924 (.a(n_3591), .b(n_2025), .y(n_3592));
nand2 g132 (.a(n_3963), .b(add_88_69_n_1530), .y(n_3591));
nor2 g131 (.a(n_3594), .b(add_88_69_n_1367), .y(n_3595));
nand2 g134 (.a(n_3593), .b(add_88_69_n_1530), .y(n_3594));
inv g135 (.a(add_88_69_n_1465), .y(n_3593));
inv g129 (.a(n_3599), .y(n_3600));
nor2 g130 (.a(n_3598), .b(n_3963), .y(n_3599));
nor2 g133 (.a(add_88_69_n_1367), .b(add_88_69_n_1465), .y(n_3598));
xor2 g209 (.a(n_3914), .b(n_3687), .y(n_3607));
nand2 g7925 (.a(n_3612), .b(n_3618), .y(n_3619));
nand2 g7926 (.a(n_3609), .b(n_3611), .y(n_3612));
nor2 g7927 (.a(n_3687), .b(n_2511), .y(n_3609));
nand2 g7929 (.a(n_3952), .b(n_3936), .y(n_3611));
nand2 g7931 (.a(n_3615), .b(n_3949), .y(n_3618));
nor2 g7932 (.a(n_3687), .b(n_3614), .y(n_3615));
inv g7933 (.a(n_3613), .y(n_3614));
nor2 g7934 (.a(n_3951), .b(n_3713), .y(n_3613));
inv g7936 (.a(n_3936), .y(n_3616));
nand2 g7937 (.a(n_3624), .b(n_1820), .y(n_3625));
nor2 g7938 (.a(n_3970), .b(n_1813), .y(n_3624));
nand2 g7943 (.a(n_3631), .b(n_3636), .y(n_3637));
nand2 g7944 (.a(n_3629), .b(n_3630), .y(n_3631));
inv g7945 (.a(n_3628), .y(n_3629));
nand2 g7946 (.a(n_3626), .b(n_3627), .y(n_3628));
nand2 g637 (.a(n_2103), .b(add_88_69_n_1456), .y(n_3626));
nor2 g634 (.a(add_88_69_n_1377), .b(v1_23_), .y(n_3627));
nor2 g636 (.a(add_88_69_n_1363), .b(n_1389), .y(n_3630));
nand2 g7947 (.a(n_3633), .b(n_3635), .y(n_3636));
nand2 g631 (.a(n_3626), .b(n_3632), .y(n_3633));
nor2 g635 (.a(add_88_69_n_1363), .b(add_88_69_n_1377), .y(n_3632));
nor2 g638 (.a(n_3634), .b(v1_23_), .y(n_3635));
inv g639 (.a(n_1389), .y(n_3634));
xor2 g7948 (.a(n_3633), .b(n_1389), .y(n_3638));
nand2 g156 (.a(n_3641), .b(n_3644), .y(n_3645));
nor2 g158 (.a(n_3640), .b(add_76_82_n_948), .y(n_3641));
nor2 g162 (.a(n_2363), .b(add_76_82_n_1070), .y(n_3640));
nand2 g159 (.a(n_3904), .b(n_3643), .y(n_3644));
nor2 g160 (.a(add_76_82_n_1070), .b(n_2798), .y(n_3643));
inv g155 (.a(n_3645), .y(n_3646));
nor2 g154 (.a(n_3648), .b(add_76_82_n_1070), .y(n_3649));
nor2 g157 (.a(n_3906), .b(add_76_82_n_954), .y(n_3648));
nor2 g56 (.a(n_3649), .b(n_3650), .y(n_3651));
inv g7951 (.a(n_2347), .y(n_3650));
xor2 g7952 (.a(n_2733), .b(n_1490), .y(n_3652));
nand2 g7953 (.a(n_3656), .b(n_3659), .y(n_3660));
nor2 g101 (.a(n_1980), .b(n_3655), .y(n_3656));
nor2 g105 (.a(add_76_21_n_1002), .b(add_76_21_n_1019), .y(n_3655));
nand2 g7954 (.a(n_3658), .b(n_2017), .y(n_3659));
nor2 g7955 (.a(add_76_21_n_1002), .b(n_3657), .y(n_3658));
inv g7956 (.a(n_2020), .y(n_3657));
nor2 g7957 (.a(n_3663), .b(add_76_21_n_1002), .y(n_3664));
inv g7958 (.a(n_3662), .y(n_3663));
nand2 g7959 (.a(n_3661), .b(add_76_21_n_1019), .y(n_3662));
nand2 g106 (.a(n_2017), .b(n_2020), .y(n_3661));
nand2 g7962 (.a(n_3667), .b(n_1895), .y(n_3668));
nand2 g39 (.a(n_3709), .b(n_1892), .y(n_3667));
nand2 g138 (.a(n_2019), .b(n_2018), .y(n_3671));
nand2 g7967 (.a(n_3678), .b(n_2019), .y(n_3679));
inv g136 (.a(n_3677), .y(n_3678));
nor2 g137 (.a(n_2018), .b(n_3694), .y(n_3677));
xor2 g7971 (.a(n_2005), .b(n_2085), .y(n_3680));
nor2 g7972 (.a(add_76_21_n_818), .b(add_76_21_n_914), .y(n_3681));
xor2 g7975 (.a(n_3681), .b(n_2085), .y(n_3687));
nand2 g7976 (.a(n_3692), .b(n_3699), .y(n_3700));
nor2 g7977 (.a(n_3689), .b(n_3691), .y(n_3692));
nor2 g7978 (.a(n_3688), .b(v0_10_), .y(n_3689));
xor2 g7979 (.a(n_1498), .b(n_3440), .y(n_3688));
nand2 g460 (.a(n_3690), .b(n_2346), .y(n_3691));
nand2 g7980 (.a(n_3651), .b(n_3652), .y(n_3690));
nor2 g7981 (.a(n_3694), .b(n_4092), .y(n_3699));
nor2 g7982 (.a(n_3693), .b(v0_9_), .y(n_3694));
xor2 g7983 (.a(n_1504), .b(n_2370), .y(n_3693));
xor2 g7986 (.a(n_2373), .b(n_3648), .y(n_3701));
xor2 g533 (.a(n_3705), .b(n_3706), .y(n_3707));
nor2 g535 (.a(n_3702), .b(n_3704), .y(n_3705));
nand2 g539 (.a(n_2743), .b(add_76_21_n_1040), .y(n_3702));
inv g537 (.a(n_3703), .y(n_3704));
nand2 g538 (.a(n_3662), .b(add_76_21_n_1068), .y(n_3703));
xor2 g536 (.a(n_3139), .b(add_76_21_n_1134), .y(n_3706));
xor2 g534 (.a(n_3705), .b(add_76_21_n_1134), .y(n_3708));
xor2 g7987 (.a(n_3710), .b(n_3711), .y(n_3712));
nor2 g7988 (.a(n_3709), .b(n_3664), .y(n_3710));
nand2 g7989 (.a(add_76_21_n_928), .b(n_2963), .y(n_3709));
xor2 g7990 (.a(n_1240), .b(add_76_21_n_1156), .y(n_3711));
xor2 g7991 (.a(n_3710), .b(add_76_21_n_1156), .y(n_3713));
nand2 g7992 (.a(n_3718), .b(n_3725), .y(n_3726));
nand2 g7993 (.a(n_3716), .b(n_3717), .y(n_3718));
inv g7994 (.a(n_3715), .y(n_3716));
nor2 g7995 (.a(n_3714), .b(add_88_69_n_1271), .y(n_3715));
nand2 g7996 (.a(add_88_69_n_1341), .b(n_3956), .y(n_3714));
nor2 g7997 (.a(n_1580), .b(v1_22_), .y(n_3717));
nand2 g7998 (.a(n_3720), .b(n_3724), .y(n_3725));
nor2 g7999 (.a(add_88_69_n_1271), .b(n_3719), .y(n_3720));
inv g8000 (.a(add_88_69_n_1341), .y(n_3719));
nor2 g8001 (.a(n_3721), .b(n_3723), .y(n_3724));
inv g8002 (.a(n_1580), .y(n_3721));
nand2 g8003 (.a(n_3956), .b(n_3722), .y(n_3723));
inv g8004 (.a(v1_22_), .y(n_3722));
xor2 g8005 (.a(n_3715), .b(n_1580), .y(n_3727));
nand2 g8006 (.a(n_3729), .b(n_3732), .y(n_3733));
nor2 g8007 (.a(n_3728), .b(add_76_21_n_890), .y(n_3729));
inv g8008 (.a(n_2832), .y(n_3728));
inv g8009 (.a(n_3731), .y(n_3732));
nor2 g8010 (.a(n_3941), .b(add_76_21_n_978), .y(n_3731));
nand2 g598 (.a(n_3737), .b(n_3743), .y(n_3744));
mux2 g8012 (.a(n_3735), .b(n_3751), .sel(n_3804), .y(n_3737));
nor2 g612 (.a(n_3734), .b(sum_12_), .y(n_3735));
nor2 g8013 (.a(n_4138), .b(n_3742), .y(n_3743));
inv g614 (.a(inc_add_77_23_n_508), .y(n_3738));
nand2 g605 (.a(n_4136), .b(key_r_64_), .y(n_3742));
nand2 g8015 (.a(n_4597), .b(n_3760), .y(n_3761));
nor2 g8020 (.a(n_3757), .b(n_3759), .y(n_3760));
nand2 g8024 (.a(n_3758), .b(key_r_32_), .y(n_3759));
nand2 g8025 (.a(inc_add_77_23_n_493), .b(n_3751), .y(n_3758));
inv g8027 (.a(n_3814), .y(n_3764));
nand2 g8032 (.a(n_3771), .b(n_3778), .y(n_3779));
inv g8033 (.a(n_3770), .y(n_3771));
mux2 g8034 (.a(n_3768), .b(n_3751), .sel(n_3804), .y(n_3770));
nand2 g692 (.a(sum_12_), .b(sum_11_), .y(n_3768));
nor2 g8035 (.a(n_4138), .b(n_3777), .y(n_3778));
nand2 g685 (.a(n_4136), .b(key_r_0_), .y(n_3777));
nand2 g8040 (.a(n_4597), .b(n_3795), .y(n_3796));
nor2 g8043 (.a(n_3792), .b(n_3794), .y(n_3795));
inv g604 (.a(n_3791), .y(n_3792));
nand2 g8044 (.a(inc_add_77_23_n_465), .b(n_3790), .y(n_3791));
nor2 g608 (.a(inc_add_77_23_n_493), .b(sum_12_), .y(n_3790));
nand2 g603 (.a(n_4055), .b(key_r_96_), .y(n_3794));
nor2 g8057 (.a(n_3804), .b(inc_add_77_23_n_508), .y(n_3805));
nand2 g8058 (.a(inc_add_77_23_n_496), .b(inc_add_77_23_n_494), .y(n_3804));
nand2 g8059 (.a(n_3973), .b(n_3813), .y(n_3814));
nand2 g8064 (.a(n_3804), .b(sum_12_), .y(n_3813));
mux2 g8066 (.a(n_3817), .b(n_3819), .sel(n_3838), .y(n_3821));
nor2 g8067 (.a(n_3814), .b(n_3816), .y(n_3817));
inv g8068 (.a(key_r_65_), .y(n_3816));
nor2 g8069 (.a(n_3764), .b(n_3818), .y(n_3819));
inv g8070 (.a(key_r_33_), .y(n_3818));
mux2 g8075 (.a(n_3826), .b(n_3828), .sel(n_3838), .y(n_3830));
inv g152 (.a(n_3825), .y(n_3826));
nand2 g153 (.a(n_3814), .b(key_r_1_), .y(n_3825));
nor2 g8076 (.a(n_3814), .b(n_3827), .y(n_3828));
inv g8077 (.a(key_r_97_), .y(n_3827));
inv g8078 (.a(n_3831), .y(n_3832));
nand2 g8079 (.a(n_3838), .b(n_3814), .y(n_3831));
nor2 g150 (.a(n_3838), .b(n_3814), .y(n_3833));
mux2 g8080 (.a(n_3835), .b(n_3837), .sel(n_3838), .y(n_3839));
nor2 g8081 (.a(n_3814), .b(n_3834), .y(n_3835));
inv g8082 (.a(key_r_66_), .y(n_3834));
nor2 g8083 (.a(n_3764), .b(n_3836), .y(n_3837));
inv g8084 (.a(key_r_34_), .y(n_3836));
xor2 g8085 (.a(n_3805), .b(sum_11_), .y(n_3838));
nor2 g8086 (.a(n_3840), .b(n_3814), .y(n_3841));
inv g8087 (.a(n_3838), .y(n_3840));
nor2 g8088 (.a(n_3838), .b(n_3764), .y(n_3842));
nor2 g8089 (.a(n_3845), .b(n_3848), .y(n_3849));
nor2 g8090 (.a(n_3843), .b(n_3844), .y(n_3845));
nand2 g8091 (.a(n_2565), .b(n_2566), .y(n_3843));
nand2 g8092 (.a(n_1647), .b(add_76_69_n_835), .y(n_3844));
mux2 g8093 (.a(n_3847), .b(add_76_69_n_836), .sel(n_1647), .y(n_3848));
nor2 g8094 (.a(add_76_69_n_836), .b(add_76_69_n_896), .y(n_3847));
inv g8095 (.a(add_76_69_n_835), .y(add_76_69_n_836));
nor2 g8096 (.a(n_3852), .b(n_3853), .y(n_3854));
nor2 g8097 (.a(n_2565), .b(n_3851), .y(n_3852));
nand2 g8098 (.a(n_3850), .b(add_76_69_n_896), .y(n_3851));
inv g8099 (.a(n_1647), .y(n_3850));
nor2 g8100 (.a(n_2566), .b(n_3851), .y(n_3853));
nor2 g201 (.a(n_2563), .b(n_4499), .y(n_3861));
nand2 g8107 (.a(n_2619), .b(add_76_82_n_896), .y(n_3866));
xor2 g8108 (.a(n_3866), .b(n_2569), .y(n_3869));
nand2 g8109 (.a(n_3874), .b(n_3880), .y(n_3881));
nand2 g8110 (.a(n_3871), .b(n_4259), .y(n_3874));
nor2 g8111 (.a(n_4258), .b(v0_18_), .y(n_3871));
nor2 g8114 (.a(n_2531), .b(add_76_82_n_1062), .y(n_3872));
nand2 g8115 (.a(n_3876), .b(n_3879), .y(n_3880));
nor2 g8116 (.a(n_4257), .b(n_3875), .y(n_3876));
inv g8117 (.a(n_2536), .y(n_3875));
nor2 g8118 (.a(n_2531), .b(n_3878), .y(n_3879));
inv g8119 (.a(n_3877), .y(n_3878));
nor2 g8120 (.a(add_76_82_n_1062), .b(v0_18_), .y(n_3877));
nor2 g8121 (.a(add_88_69_n_1632), .b(n_3886), .y(n_3887));
nor2 g8122 (.a(n_4303), .b(n_3454), .y(n_3886));
xor2 g8126 (.a(n_4306), .b(n_1235), .y(n_3888));
nor2 g8127 (.a(n_3890), .b(n_3893), .y(n_3894));
nand2 g44 (.a(add_88_21_n_693), .b(n_2846), .y(n_3890));
inv g8129 (.a(n_3892), .y(n_3893));
nor2 g8130 (.a(n_3891), .b(n_4031), .y(n_3892));
nand2 g43 (.a(add_88_21_n_917), .b(add_88_21_n_929), .y(n_3891));
inv g218 (.a(n_3900), .y(n_3901));
nor2 g219 (.a(n_3968), .b(n_3964), .y(n_3900));
nand2 g8132 (.a(n_2842), .b(n_3895), .y(n_3896));
inv g8133 (.a(add_88_69_n_1739), .y(n_3895));
nor2 g8135 (.a(n_3905), .b(n_2798), .y(n_3906));
inv g166 (.a(n_3904), .y(n_3905));
nand2 g167 (.a(n_3902), .b(n_3903), .y(n_3904));
nand2 g168 (.a(n_4350), .b(n_2915), .y(n_3902));
nand2 g169 (.a(n_2903), .b(n_2905), .y(n_3903));
nor2 g8136 (.a(n_3905), .b(n_2356), .y(n_3907));
nor2 g8137 (.a(n_2576), .b(n_3905), .y(n_3908));
nand2 g8138 (.a(n_3904), .b(n_2805), .y(n_3909));
nand2 g8139 (.a(n_3904), .b(add_76_82_n_1066), .y(n_3910));
nand2 g8140 (.a(n_3904), .b(add_76_82_n_1088), .y(n_3911));
nand2 g8141 (.a(n_3902), .b(n_2696), .y(n_3912));
nand2 g165 (.a(n_3903), .b(add_76_82_n_1144), .y(n_3913));
xor2 g8142 (.a(n_2675), .b(add_76_21_n_1155), .y(n_3914));
nor2 g8150 (.a(n_4062), .b(n_2096), .y(n_3926));
nand2 g140 (.a(add_76_21_n_963), .b(add_76_21_n_1047), .y(n_3927));
nor2 g142 (.a(add_76_21_n_1003), .b(add_76_21_n_915), .y(n_3928));
nor2 g8152 (.a(n_1941), .b(n_3935), .y(n_3936));
nor2 g8153 (.a(n_3932), .b(n_3934), .y(n_3935));
nand2 g8154 (.a(n_3931), .b(add_76_21_n_963), .y(n_3932));
inv g8155 (.a(n_3930), .y(n_3931));
nand2 g8156 (.a(add_76_21_n_1047), .b(n_1935), .y(n_3930));
nand2 g139 (.a(add_76_21_n_950), .b(n_3933), .y(n_3934));
inv g141 (.a(n_3928), .y(n_3933));
nor2 g362 (.a(n_3927), .b(n_3928), .y(n_3941));
nor2 g8161 (.a(n_3616), .b(n_3948), .y(n_3949));
nand2 g8162 (.a(n_3946), .b(n_3947), .y(n_3948));
inv g8163 (.a(n_3945), .y(n_3946));
nand2 g8164 (.a(n_3943), .b(n_3944), .y(n_3945));
nand2 g8165 (.a(n_3928), .b(n_3942), .y(n_3943));
nor2 g8166 (.a(n_1924), .b(n_1605), .y(n_3942));
nor2 g363 (.a(n_1930), .b(n_1931), .y(n_3944));
nand2 g8167 (.a(n_3927), .b(n_3942), .y(n_3947));
nor2 g8168 (.a(n_3951), .b(n_3948), .y(n_3952));
nor2 g8169 (.a(n_1936), .b(n_3950), .y(n_3951));
inv g8170 (.a(n_3941), .y(n_3950));
inv g8171 (.a(n_3948), .y(n_3953));
nor2 g8172 (.a(n_1959), .b(n_3950), .y(n_3954));
nand2 g8173 (.a(add_76_21_n_949), .b(n_3942), .y(n_3955));
nor2 g8174 (.a(n_2204), .b(n_4062), .y(n_3956));
nand2 g8175 (.a(add_88_69_n_1341), .b(n_3961), .y(n_3962));
nor2 g8176 (.a(n_3958), .b(n_3960), .y(n_3961));
nand2 g8177 (.a(n_3956), .b(n_4100), .y(n_3958));
inv g8179 (.a(n_3959), .y(n_3960));
nor2 g8180 (.a(n_3575), .b(add_88_69_n_1634), .y(n_3959));
nand2 g8181 (.a(add_88_69_n_1424), .b(n_3959), .y(n_3963));
nor2 g8182 (.a(n_3959), .b(add_88_69_n_1739), .y(n_3964));
nor2 g8183 (.a(add_88_69_n_1739), .b(n_3965), .y(n_3966));
inv g8184 (.a(n_4100), .y(n_3965));
nor2 g8185 (.a(add_88_69_n_1647), .b(n_4100), .y(n_3967));
nand2 g8186 (.a(n_3896), .b(n_4100), .y(n_3968));
nor2 g8187 (.a(n_3969), .b(n_1810), .y(n_3970));
nand2 g8188 (.a(n_1808), .b(add_88_21_n_688), .y(n_3969));
inv g4 (.a(n_3972), .y(n_3973));
nand2 g8189 (.a(n_4055), .b(n_3791), .y(n_3972));
nand2 g8191 (.a(n_3974), .b(add_88_82_n_1967), .y(n_3975));
nor2 g8192 (.a(add_88_82_n_2288), .b(add_88_82_n_2042), .y(n_3974));
nand2 add_88_82_g8193 (.a(add_88_82_n_1967), .b(n_3976), .y(n_3977));
inv add_88_82_g8194 (.a(add_88_82_n_2288), .y(n_3976));
xor2 g6402__8195 (.a(n_3982), .b(n_3008), .y(n_3983));
xor2 add_76_82_g8196 (.a(n_3980), .b(n_3981), .y(n_3982));
xor2 add_76_69_g8197 (.a(n_3978), .b(n_3979), .y(n_3980));
nor2 add_76_82_g8198 (.a(add_76_82_n_1218), .b(add_76_82_n_1296), .y(n_3978));
nor2 add_76_69_g8199 (.a(add_76_69_n_1099), .b(add_76_69_n_1105), .y(n_3979));
nand2 add_76_69_g8200 (.a(add_76_69_n_669), .b(add_76_69_n_661), .y(n_3981));
nor2 g8201 (.a(add_76_82_n_840), .b(add_76_82_n_855), .y(n_3984));
nand2 g8202 (.a(add_76_82_n_1259), .b(add_76_82_n_1213), .y(n_3985));
xor2 g8203 (.a(n_2044), .b(n_2045), .y(n_3986));
nand2 add_76_21_g8204 (.a(n_3988), .b(v0_29_), .y(n_3989));
xor2 g8205 (.a(n_4058), .b(n_3984), .y(n_3988));
nor2 g8214 (.a(n_4001), .b(n_4371), .y(n_4002));
xor2 g8215 (.a(n_3997), .b(n_4000), .y(n_4001));
nand2 add_88_69_g1548__8216 (.a(add_88_69_n_1289), .b(add_88_69_n_1267), .y(n_3997));
xor2 add_88_69_g1539__8217 (.a(n_3998), .b(n_3999), .y(n_4000));
xor2 g8218 (.a(n_2982), .b(n_2983), .y(n_3998));
xor2 add_88_69_g8219 (.a(n_1216), .b(n_3525), .y(n_3999));
nand2 g8220 (.a(n_4001), .b(n_1683), .y(n_4003));
nand2 g8234 (.a(n_4025), .b(n_4030), .y(n_4031));
nand2 g8235 (.a(n_4019), .b(n_4024), .y(n_4025));
nand2 g619 (.a(n_4017), .b(n_4018), .y(n_4019));
nor2 g8236 (.a(add_88_69_n_1315), .b(n_1919), .y(n_4017));
nand2 g8237 (.a(add_88_69_n_1395), .b(n_2103), .y(n_4018));
nor2 g616 (.a(n_4023), .b(v1_28_), .y(n_4024));
inv g617 (.a(n_4022), .y(n_4023));
xor2 g618 (.a(n_4020), .b(n_4021), .y(n_4022));
xor2 g622 (.a(add_88_82_n_1906), .b(add_88_82_n_2142), .y(n_4020));
nor2 g8238 (.a(n_1904), .b(n_2035), .y(n_4021));
nand2 g8239 (.a(n_4028), .b(n_4029), .y(n_4030));
inv g620 (.a(n_4027), .y(n_4028));
nand2 g621 (.a(n_4026), .b(n_4018), .y(n_4027));
nor2 g624 (.a(n_1919), .b(v1_28_), .y(n_4026));
nor2 g615 (.a(add_88_69_n_1315), .b(n_4022), .y(n_4029));
inv g8254 (.a(n_3571), .y(n_4048));
nor2 g8255 (.a(n_4046), .b(n_3668), .y(n_3571));
nand2 g8256 (.a(n_3527), .b(n_1890), .y(n_4046));
inv g8257 (.a(n_3527), .y(n_4049));
nand2 g8263 (.a(inc_add_77_23_n_493), .b(sum_12_), .y(n_4055));
xor2 g8265 (.a(inc_add_77_23_n_508), .b(sum_11_), .y(n_4057));
xor2 g8266 (.a(n_3986), .b(n_3985), .y(n_4058));
xor2 g8267 (.a(n_3490), .b(n_3491), .y(n_4059));
inv g8268 (.a(n_4061), .y(n_4062));
nand2 g8269 (.a(n_4060), .b(n_4306), .y(n_4061));
xor2 g8270 (.a(n_4059), .b(n_3493), .y(n_4060));
nor2 g8295 (.a(n_4087), .b(n_3505), .y(n_4088));
xor2 g8296 (.a(n_3520), .b(n_3514), .y(n_4087));
nand2 g8297 (.a(n_4089), .b(n_1998), .y(n_4090));
xor2 g8298 (.a(n_3680), .b(n_3681), .y(n_4089));
nor2 g8299 (.a(n_4091), .b(v0_8_), .y(n_4092));
mux2 g8300 (.a(n_2362), .b(n_3648), .sel(n_2373), .y(n_4091));
nand2 g8307 (.a(n_4099), .b(n_2033), .y(n_4100));
mux2 g8308 (.a(n_2517), .b(n_3687), .sel(n_3914), .y(n_4099));
nand2 inc_add_77_23_g8342 (.a(inc_add_77_23_n_492), .b(sum_12_), .y(n_4135));
nand2 g8343 (.a(inc_add_77_23_n_508), .b(n_3734), .y(n_4136));
nand2 g8344 (.a(n_3738), .b(sum_11_), .y(n_4137));
nor2 g8345 (.a(n_3804), .b(n_4137), .y(n_4138));
inv g8403 (.a(sum_12_), .y(n_3751));
inv g8404 (.a(sum_11_), .y(n_3734));
inv g8407 (.a(n_4135), .y(n_3757));
inv g8470 (.a(n_4257), .y(n_4258));
nand2 g8471 (.a(n_3849), .b(n_3854), .y(n_4257));
nand2 g8472 (.a(n_3872), .b(n_2536), .y(n_4259));
inv g839 (.a(n_4289), .y(n_4290));
nor2 g840 (.a(n_4283), .b(n_4502), .y(n_4289));
nor2 g8489 (.a(n_4279), .b(n_4282), .y(n_4283));
nand2 g842 (.a(n_4277), .b(n_4278), .y(n_4279));
xor2 g847 (.a(n_3866), .b(n_2569), .y(n_4277));
nand2 g848 (.a(n_2771), .b(n_2772), .y(n_4278));
nand2 g845 (.a(n_4281), .b(v0_16_), .y(n_4282));
inv g851 (.a(n_4280), .y(n_4281));
nor2 g852 (.a(n_2766), .b(n_2761), .y(n_4280));
nand2 g846 (.a(n_4281), .b(n_4278), .y(n_4291));
nand2 g8493 (.a(n_4277), .b(v0_16_), .y(n_4292));
nand2 g834 (.a(n_4298), .b(n_4302), .y(n_4303));
mux2 g835 (.a(n_4295), .b(n_4296), .sel(n_4297), .y(n_4298));
nand2 g8494 (.a(n_4293), .b(n_4294), .y(n_4295));
nor2 g8495 (.a(n_1235), .b(n_2828), .y(n_4293));
inv g8496 (.a(n_2815), .y(n_4294));
inv g8497 (.a(n_1235), .y(n_4296));
nor2 g8498 (.a(n_2821), .b(n_2825), .y(n_4297));
nor2 g836 (.a(n_4300), .b(n_4301), .y(n_4302));
nand2 g838 (.a(n_3713), .b(n_4299), .y(n_4300));
nand2 g8499 (.a(n_1235), .b(n_2828), .y(n_4299));
nor2 g8500 (.a(n_4294), .b(n_4296), .y(n_4301));
nand2 g837 (.a(n_4304), .b(n_4305), .y(n_4306));
nor2 g8501 (.a(n_2821), .b(n_2815), .y(n_4304));
nor2 g8502 (.a(n_2825), .b(n_2828), .y(n_4305));
nand2 g8526 (.a(n_4335), .b(n_4336), .y(n_4337));
mux2 g8527 (.a(n_4332), .b(n_4334), .sel(add_88_21_n_812), .y(n_4335));
inv g8528 (.a(n_4331), .y(n_4332));
nor2 g8529 (.a(add_88_21_n_982), .b(n_4371), .y(n_4331));
nand2 g8531 (.a(add_88_21_n_982), .b(n_1683), .y(n_4334));
nand2 g8533 (.a(n_4371), .b(v1_r_3_), .y(n_4336));
nand2 g8543 (.a(n_1870), .b(n_1861), .y(n_4350));
nor2 add_76_21_g8544 (.a(n_4354), .b(v0_2_), .y(n_4355));
xor2 g6427__8545 (.a(n_4353), .b(n_4350), .y(n_4354));
xor2 g8546 (.a(n_4351), .b(n_4352), .y(n_4353));
xor2 add_76_69_g8547 (.a(add_76_69_n_869), .b(add_76_69_n_952), .y(n_4351));
nor2 add_76_82_g8548 (.a(add_76_82_n_1287), .b(n_2681), .y(n_4352));
nand2 add_76_21_g8549 (.a(n_4354), .b(v0_2_), .y(n_4356));
nor2 g8553 (.a(add_88_21_n_987), .b(n_4371), .y(n_4358));
nand2 g8557 (.a(n_4371), .b(v1_r_5_), .y(n_4363));
mux2 g8558 (.a(n_4366), .b(n_4368), .sel(n_4369), .y(n_4370));
nand2 g7590_dup2 (.a(n_4365), .b(n_3177), .y(n_4366));
inv g8559 (.a(n_3172), .y(n_4365));
nand2 g8560 (.a(n_4367), .b(n_3177), .y(n_4368));
nand2 g8561 (.a(add_88_21_n_1014), .b(n_1683), .y(n_4367));
nand2 add_88_21_g8562 (.a(add_88_21_n_900), .b(add_88_21_n_753), .y(n_4369));
nor2 g8566 (.a(add_88_21_n_1013), .b(n_4371), .y(n_4372));
nand2 g8567 (.a(ps_1_), .b(n_1800), .y(n_4371));
nand2 g93 (.a(n_4371), .b(v1_r_7_), .y(n_4377));
nand2 g8572 (.a(add_88_21_n_830), .b(add_88_21_n_727), .y(n_4380));
nand2 g8586 (.a(n_4397), .b(n_3671), .y(n_4398));
nor2 g8587 (.a(n_3689), .b(n_3694), .y(n_4397));
inv add_76_21_g8588 (.a(n_3689), .y(n_4399));
mux2 g8589 (.a(n_4401), .b(n_4403), .sel(n_4404), .y(n_4405));
nand2 g8550_dup2 (.a(n_4400), .b(n_4363), .y(n_4401));
inv g8590 (.a(n_4358), .y(n_4400));
nand2 g8591 (.a(n_4402), .b(n_4363), .y(n_4403));
nand2 g8592 (.a(add_88_21_n_987), .b(n_1683), .y(n_4402));
nand2 add_88_21_g8593 (.a(add_88_21_n_756), .b(add_88_21_n_1042), .y(n_4404));
mux2 g8594 (.a(n_4407), .b(n_4409), .sel(n_4410), .y(n_4411));
nand2 g8563_dup2 (.a(n_4406), .b(n_4377), .y(n_4407));
inv g8595 (.a(n_4372), .y(n_4406));
nand2 g8596 (.a(n_4408), .b(n_4377), .y(n_4409));
nand2 g8597 (.a(add_88_21_n_1013), .b(n_1683), .y(n_4408));
nor2 add_88_21_g8598 (.a(add_88_21_n_801), .b(add_88_21_n_733), .y(n_4410));
nand2 g8685 (.a(n_4498), .b(v0_18_), .y(n_4499));
mux2 g8686 (.a(n_4258), .b(n_4257), .sel(n_4259), .y(n_4498));
inv g8687 (.a(n_4501), .y(n_4502));
nand2 g8688 (.a(n_4500), .b(v0_17_), .y(n_4501));
xor2 g8689 (.a(n_2766), .b(n_2772), .y(n_4500));
nor2 g8733 (.a(n_4549), .b(add_88_21_n_772), .y(n_4550));
nand2 g8734 (.a(n_4380), .b(add_88_21_n_1053), .y(n_4549));
mux2 g8735 (.a(n_3372), .b(n_3370), .sel(n_4550), .y(n_4552));
inv g8740 (.a(n_4557), .y(n_4558));
nor2 g8741 (.a(n_1528), .b(add_76_69_n_1090), .y(n_4557));
mux2 g8780 (.a(n_3734), .b(n_4057), .sel(n_3804), .y(n_4597));
endmodule

